module RandomLUT(
  input  [11:0] io_in,
  output [11:0] io_out
);
  wire [11:0] _GEN_1 = 12'h1 == io_in ? 12'h939 : 12'hded; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2 = 12'h2 == io_in ? 12'he75 : _GEN_1; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3 = 12'h3 == io_in ? 12'h431 : _GEN_2; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4 = 12'h4 == io_in ? 12'h874 : _GEN_3; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_5 = 12'h5 == io_in ? 12'hb42 : _GEN_4; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_6 = 12'h6 == io_in ? 12'h53f : _GEN_5; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_7 = 12'h7 == io_in ? 12'h4b1 : _GEN_6; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_8 = 12'h8 == io_in ? 12'hd03 : _GEN_7; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_9 = 12'h9 == io_in ? 12'h70c : _GEN_8; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_10 = 12'ha == io_in ? 12'hf46 : _GEN_9; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_11 = 12'hb == io_in ? 12'hf41 : _GEN_10; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_12 = 12'hc == io_in ? 12'h655 : _GEN_11; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_13 = 12'hd == io_in ? 12'haa1 : _GEN_12; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_14 = 12'he == io_in ? 12'h71c : _GEN_13; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_15 = 12'hf == io_in ? 12'h863 : _GEN_14; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_16 = 12'h10 == io_in ? 12'h22e : _GEN_15; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_17 = 12'h11 == io_in ? 12'h70a : _GEN_16; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_18 = 12'h12 == io_in ? 12'hc60 : _GEN_17; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_19 = 12'h13 == io_in ? 12'hfda : _GEN_18; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_20 = 12'h14 == io_in ? 12'h3de : _GEN_19; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_21 = 12'h15 == io_in ? 12'h38c : _GEN_20; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_22 = 12'h16 == io_in ? 12'haa2 : _GEN_21; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_23 = 12'h17 == io_in ? 12'h8ea : _GEN_22; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_24 = 12'h18 == io_in ? 12'h9b2 : _GEN_23; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_25 = 12'h19 == io_in ? 12'hc34 : _GEN_24; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_26 = 12'h1a == io_in ? 12'h31 : _GEN_25; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_27 = 12'h1b == io_in ? 12'h5d5 : _GEN_26; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_28 = 12'h1c == io_in ? 12'h431 : _GEN_27; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_29 = 12'h1d == io_in ? 12'h2d : _GEN_28; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_30 = 12'h1e == io_in ? 12'hfb0 : _GEN_29; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_31 = 12'h1f == io_in ? 12'he5e : _GEN_30; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_32 = 12'h20 == io_in ? 12'h7c8 : _GEN_31; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_33 = 12'h21 == io_in ? 12'hd5f : _GEN_32; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_34 = 12'h22 == io_in ? 12'h46 : _GEN_33; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_35 = 12'h23 == io_in ? 12'hb18 : _GEN_34; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_36 = 12'h24 == io_in ? 12'he86 : _GEN_35; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_37 = 12'h25 == io_in ? 12'h7c4 : _GEN_36; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_38 = 12'h26 == io_in ? 12'h9fb : _GEN_37; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_39 = 12'h27 == io_in ? 12'h342 : _GEN_38; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_40 = 12'h28 == io_in ? 12'ha33 : _GEN_39; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_41 = 12'h29 == io_in ? 12'ha3e : _GEN_40; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_42 = 12'h2a == io_in ? 12'h144 : _GEN_41; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_43 = 12'h2b == io_in ? 12'h248 : _GEN_42; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_44 = 12'h2c == io_in ? 12'h1aa : _GEN_43; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_45 = 12'h2d == io_in ? 12'h966 : _GEN_44; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_46 = 12'h2e == io_in ? 12'hbd5 : _GEN_45; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_47 = 12'h2f == io_in ? 12'h635 : _GEN_46; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_48 = 12'h30 == io_in ? 12'hbda : _GEN_47; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_49 = 12'h31 == io_in ? 12'hdda : _GEN_48; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_50 = 12'h32 == io_in ? 12'h319 : _GEN_49; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_51 = 12'h33 == io_in ? 12'hf56 : _GEN_50; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_52 = 12'h34 == io_in ? 12'hbaa : _GEN_51; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_53 = 12'h35 == io_in ? 12'hca : _GEN_52; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_54 = 12'h36 == io_in ? 12'ha5b : _GEN_53; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_55 = 12'h37 == io_in ? 12'h8be : _GEN_54; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_56 = 12'h38 == io_in ? 12'ha4a : _GEN_55; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_57 = 12'h39 == io_in ? 12'h9d6 : _GEN_56; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_58 = 12'h3a == io_in ? 12'h17 : _GEN_57; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_59 = 12'h3b == io_in ? 12'h3d1 : _GEN_58; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_60 = 12'h3c == io_in ? 12'h758 : _GEN_59; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_61 = 12'h3d == io_in ? 12'hf65 : _GEN_60; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_62 = 12'h3e == io_in ? 12'h5a0 : _GEN_61; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_63 = 12'h3f == io_in ? 12'hfc : _GEN_62; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_64 = 12'h40 == io_in ? 12'h30c : _GEN_63; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_65 = 12'h41 == io_in ? 12'h1fb : _GEN_64; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_66 = 12'h42 == io_in ? 12'hd01 : _GEN_65; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_67 = 12'h43 == io_in ? 12'hba9 : _GEN_66; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_68 = 12'h44 == io_in ? 12'h693 : _GEN_67; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_69 = 12'h45 == io_in ? 12'he9b : _GEN_68; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_70 = 12'h46 == io_in ? 12'h406 : _GEN_69; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_71 = 12'h47 == io_in ? 12'hef5 : _GEN_70; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_72 = 12'h48 == io_in ? 12'h780 : _GEN_71; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_73 = 12'h49 == io_in ? 12'hc13 : _GEN_72; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_74 = 12'h4a == io_in ? 12'h1f5 : _GEN_73; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_75 = 12'h4b == io_in ? 12'he6c : _GEN_74; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_76 = 12'h4c == io_in ? 12'h66 : _GEN_75; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_77 = 12'h4d == io_in ? 12'h2a1 : _GEN_76; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_78 = 12'h4e == io_in ? 12'h2e5 : _GEN_77; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_79 = 12'h4f == io_in ? 12'hdd3 : _GEN_78; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_80 = 12'h50 == io_in ? 12'h121 : _GEN_79; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_81 = 12'h51 == io_in ? 12'h566 : _GEN_80; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_82 = 12'h52 == io_in ? 12'h462 : _GEN_81; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_83 = 12'h53 == io_in ? 12'h4ab : _GEN_82; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_84 = 12'h54 == io_in ? 12'h44f : _GEN_83; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_85 = 12'h55 == io_in ? 12'h105 : _GEN_84; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_86 = 12'h56 == io_in ? 12'h71 : _GEN_85; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_87 = 12'h57 == io_in ? 12'hd5f : _GEN_86; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_88 = 12'h58 == io_in ? 12'hdc6 : _GEN_87; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_89 = 12'h59 == io_in ? 12'hcaf : _GEN_88; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_90 = 12'h5a == io_in ? 12'h105 : _GEN_89; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_91 = 12'h5b == io_in ? 12'h184 : _GEN_90; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_92 = 12'h5c == io_in ? 12'h925 : _GEN_91; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_93 = 12'h5d == io_in ? 12'h1ce : _GEN_92; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_94 = 12'h5e == io_in ? 12'h29c : _GEN_93; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_95 = 12'h5f == io_in ? 12'h7d : _GEN_94; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_96 = 12'h60 == io_in ? 12'hbb6 : _GEN_95; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_97 = 12'h61 == io_in ? 12'hd92 : _GEN_96; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_98 = 12'h62 == io_in ? 12'h263 : _GEN_97; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_99 = 12'h63 == io_in ? 12'h51f : _GEN_98; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_100 = 12'h64 == io_in ? 12'hd63 : _GEN_99; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_101 = 12'h65 == io_in ? 12'he70 : _GEN_100; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_102 = 12'h66 == io_in ? 12'hd86 : _GEN_101; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_103 = 12'h67 == io_in ? 12'ha98 : _GEN_102; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_104 = 12'h68 == io_in ? 12'hff8 : _GEN_103; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_105 = 12'h69 == io_in ? 12'h93b : _GEN_104; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_106 = 12'h6a == io_in ? 12'h3d2 : _GEN_105; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_107 = 12'h6b == io_in ? 12'h61d : _GEN_106; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_108 = 12'h6c == io_in ? 12'h8ac : _GEN_107; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_109 = 12'h6d == io_in ? 12'h6cd : _GEN_108; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_110 = 12'h6e == io_in ? 12'h8f8 : _GEN_109; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_111 = 12'h6f == io_in ? 12'hf37 : _GEN_110; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_112 = 12'h70 == io_in ? 12'h6a4 : _GEN_111; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_113 = 12'h71 == io_in ? 12'h6fc : _GEN_112; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_114 = 12'h72 == io_in ? 12'hbac : _GEN_113; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_115 = 12'h73 == io_in ? 12'hdcb : _GEN_114; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_116 = 12'h74 == io_in ? 12'h2b8 : _GEN_115; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_117 = 12'h75 == io_in ? 12'h1c6 : _GEN_116; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_118 = 12'h76 == io_in ? 12'h1 : _GEN_117; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_119 = 12'h77 == io_in ? 12'hd36 : _GEN_118; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_120 = 12'h78 == io_in ? 12'h49c : _GEN_119; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_121 = 12'h79 == io_in ? 12'h751 : _GEN_120; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_122 = 12'h7a == io_in ? 12'h7f9 : _GEN_121; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_123 = 12'h7b == io_in ? 12'h517 : _GEN_122; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_124 = 12'h7c == io_in ? 12'h2eb : _GEN_123; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_125 = 12'h7d == io_in ? 12'h4d8 : _GEN_124; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_126 = 12'h7e == io_in ? 12'hffb : _GEN_125; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_127 = 12'h7f == io_in ? 12'h16c : _GEN_126; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_128 = 12'h80 == io_in ? 12'hc34 : _GEN_127; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_129 = 12'h81 == io_in ? 12'h3e7 : _GEN_128; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_130 = 12'h82 == io_in ? 12'h39 : _GEN_129; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_131 = 12'h83 == io_in ? 12'h738 : _GEN_130; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_132 = 12'h84 == io_in ? 12'h523 : _GEN_131; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_133 = 12'h85 == io_in ? 12'hc98 : _GEN_132; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_134 = 12'h86 == io_in ? 12'h4aa : _GEN_133; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_135 = 12'h87 == io_in ? 12'hbb8 : _GEN_134; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_136 = 12'h88 == io_in ? 12'h32e : _GEN_135; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_137 = 12'h89 == io_in ? 12'h7e1 : _GEN_136; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_138 = 12'h8a == io_in ? 12'hcd7 : _GEN_137; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_139 = 12'h8b == io_in ? 12'ha03 : _GEN_138; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_140 = 12'h8c == io_in ? 12'h476 : _GEN_139; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_141 = 12'h8d == io_in ? 12'h6d6 : _GEN_140; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_142 = 12'h8e == io_in ? 12'h656 : _GEN_141; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_143 = 12'h8f == io_in ? 12'hcc7 : _GEN_142; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_144 = 12'h90 == io_in ? 12'h784 : _GEN_143; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_145 = 12'h91 == io_in ? 12'hcb5 : _GEN_144; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_146 = 12'h92 == io_in ? 12'h90e : _GEN_145; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_147 = 12'h93 == io_in ? 12'hbd5 : _GEN_146; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_148 = 12'h94 == io_in ? 12'haca : _GEN_147; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_149 = 12'h95 == io_in ? 12'he74 : _GEN_148; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_150 = 12'h96 == io_in ? 12'h451 : _GEN_149; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_151 = 12'h97 == io_in ? 12'hb1f : _GEN_150; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_152 = 12'h98 == io_in ? 12'h233 : _GEN_151; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_153 = 12'h99 == io_in ? 12'h9a4 : _GEN_152; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_154 = 12'h9a == io_in ? 12'hef6 : _GEN_153; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_155 = 12'h9b == io_in ? 12'hb36 : _GEN_154; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_156 = 12'h9c == io_in ? 12'hd5f : _GEN_155; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_157 = 12'h9d == io_in ? 12'h107 : _GEN_156; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_158 = 12'h9e == io_in ? 12'ha65 : _GEN_157; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_159 = 12'h9f == io_in ? 12'h23a : _GEN_158; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_160 = 12'ha0 == io_in ? 12'hb74 : _GEN_159; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_161 = 12'ha1 == io_in ? 12'h5f7 : _GEN_160; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_162 = 12'ha2 == io_in ? 12'he9e : _GEN_161; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_163 = 12'ha3 == io_in ? 12'h50d : _GEN_162; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_164 = 12'ha4 == io_in ? 12'h1be : _GEN_163; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_165 = 12'ha5 == io_in ? 12'h69d : _GEN_164; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_166 = 12'ha6 == io_in ? 12'h242 : _GEN_165; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_167 = 12'ha7 == io_in ? 12'hfca : _GEN_166; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_168 = 12'ha8 == io_in ? 12'ha86 : _GEN_167; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_169 = 12'ha9 == io_in ? 12'hc5 : _GEN_168; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_170 = 12'haa == io_in ? 12'h91d : _GEN_169; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_171 = 12'hab == io_in ? 12'h395 : _GEN_170; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_172 = 12'hac == io_in ? 12'h464 : _GEN_171; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_173 = 12'had == io_in ? 12'hcff : _GEN_172; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_174 = 12'hae == io_in ? 12'h318 : _GEN_173; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_175 = 12'haf == io_in ? 12'h88 : _GEN_174; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_176 = 12'hb0 == io_in ? 12'h456 : _GEN_175; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_177 = 12'hb1 == io_in ? 12'h435 : _GEN_176; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_178 = 12'hb2 == io_in ? 12'h6ac : _GEN_177; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_179 = 12'hb3 == io_in ? 12'h9f3 : _GEN_178; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_180 = 12'hb4 == io_in ? 12'h31d : _GEN_179; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_181 = 12'hb5 == io_in ? 12'h919 : _GEN_180; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_182 = 12'hb6 == io_in ? 12'h116 : _GEN_181; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_183 = 12'hb7 == io_in ? 12'h816 : _GEN_182; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_184 = 12'hb8 == io_in ? 12'h80d : _GEN_183; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_185 = 12'hb9 == io_in ? 12'hdcd : _GEN_184; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_186 = 12'hba == io_in ? 12'h3c3 : _GEN_185; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_187 = 12'hbb == io_in ? 12'heb1 : _GEN_186; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_188 = 12'hbc == io_in ? 12'hfcf : _GEN_187; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_189 = 12'hbd == io_in ? 12'hb18 : _GEN_188; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_190 = 12'hbe == io_in ? 12'hca0 : _GEN_189; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_191 = 12'hbf == io_in ? 12'h5ec : _GEN_190; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_192 = 12'hc0 == io_in ? 12'h6c4 : _GEN_191; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_193 = 12'hc1 == io_in ? 12'h984 : _GEN_192; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_194 = 12'hc2 == io_in ? 12'hc8b : _GEN_193; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_195 = 12'hc3 == io_in ? 12'h1f7 : _GEN_194; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_196 = 12'hc4 == io_in ? 12'he01 : _GEN_195; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_197 = 12'hc5 == io_in ? 12'h43f : _GEN_196; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_198 = 12'hc6 == io_in ? 12'hda9 : _GEN_197; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_199 = 12'hc7 == io_in ? 12'hc63 : _GEN_198; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_200 = 12'hc8 == io_in ? 12'h440 : _GEN_199; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_201 = 12'hc9 == io_in ? 12'h1ed : _GEN_200; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_202 = 12'hca == io_in ? 12'hfbd : _GEN_201; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_203 = 12'hcb == io_in ? 12'hbc9 : _GEN_202; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_204 = 12'hcc == io_in ? 12'h551 : _GEN_203; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_205 = 12'hcd == io_in ? 12'h84f : _GEN_204; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_206 = 12'hce == io_in ? 12'h29f : _GEN_205; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_207 = 12'hcf == io_in ? 12'he57 : _GEN_206; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_208 = 12'hd0 == io_in ? 12'h1e8 : _GEN_207; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_209 = 12'hd1 == io_in ? 12'hd00 : _GEN_208; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_210 = 12'hd2 == io_in ? 12'ha6d : _GEN_209; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_211 = 12'hd3 == io_in ? 12'h24b : _GEN_210; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_212 = 12'hd4 == io_in ? 12'h593 : _GEN_211; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_213 = 12'hd5 == io_in ? 12'h7b6 : _GEN_212; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_214 = 12'hd6 == io_in ? 12'h401 : _GEN_213; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_215 = 12'hd7 == io_in ? 12'h3fc : _GEN_214; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_216 = 12'hd8 == io_in ? 12'hac1 : _GEN_215; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_217 = 12'hd9 == io_in ? 12'h2a2 : _GEN_216; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_218 = 12'hda == io_in ? 12'hcf6 : _GEN_217; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_219 = 12'hdb == io_in ? 12'h33 : _GEN_218; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_220 = 12'hdc == io_in ? 12'h624 : _GEN_219; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_221 = 12'hdd == io_in ? 12'hbbb : _GEN_220; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_222 = 12'hde == io_in ? 12'h5bc : _GEN_221; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_223 = 12'hdf == io_in ? 12'hfeb : _GEN_222; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_224 = 12'he0 == io_in ? 12'hf7d : _GEN_223; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_225 = 12'he1 == io_in ? 12'h2c : _GEN_224; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_226 = 12'he2 == io_in ? 12'heb7 : _GEN_225; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_227 = 12'he3 == io_in ? 12'h85 : _GEN_226; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_228 = 12'he4 == io_in ? 12'h198 : _GEN_227; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_229 = 12'he5 == io_in ? 12'h218 : _GEN_228; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_230 = 12'he6 == io_in ? 12'h601 : _GEN_229; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_231 = 12'he7 == io_in ? 12'h283 : _GEN_230; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_232 = 12'he8 == io_in ? 12'hc5f : _GEN_231; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_233 = 12'he9 == io_in ? 12'h2e0 : _GEN_232; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_234 = 12'hea == io_in ? 12'h200 : _GEN_233; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_235 = 12'heb == io_in ? 12'h5cf : _GEN_234; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_236 = 12'hec == io_in ? 12'hc9 : _GEN_235; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_237 = 12'hed == io_in ? 12'h290 : _GEN_236; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_238 = 12'hee == io_in ? 12'he65 : _GEN_237; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_239 = 12'hef == io_in ? 12'hb38 : _GEN_238; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_240 = 12'hf0 == io_in ? 12'hfe0 : _GEN_239; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_241 = 12'hf1 == io_in ? 12'ha5a : _GEN_240; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_242 = 12'hf2 == io_in ? 12'hc04 : _GEN_241; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_243 = 12'hf3 == io_in ? 12'h8fb : _GEN_242; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_244 = 12'hf4 == io_in ? 12'h4b6 : _GEN_243; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_245 = 12'hf5 == io_in ? 12'he28 : _GEN_244; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_246 = 12'hf6 == io_in ? 12'hfa7 : _GEN_245; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_247 = 12'hf7 == io_in ? 12'h566 : _GEN_246; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_248 = 12'hf8 == io_in ? 12'h8c9 : _GEN_247; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_249 = 12'hf9 == io_in ? 12'hbb1 : _GEN_248; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_250 = 12'hfa == io_in ? 12'hd4e : _GEN_249; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_251 = 12'hfb == io_in ? 12'h601 : _GEN_250; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_252 = 12'hfc == io_in ? 12'h5b7 : _GEN_251; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_253 = 12'hfd == io_in ? 12'h5da : _GEN_252; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_254 = 12'hfe == io_in ? 12'h286 : _GEN_253; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_255 = 12'hff == io_in ? 12'h8cf : _GEN_254; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_256 = 12'h100 == io_in ? 12'h486 : _GEN_255; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_257 = 12'h101 == io_in ? 12'h616 : _GEN_256; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_258 = 12'h102 == io_in ? 12'h6c6 : _GEN_257; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_259 = 12'h103 == io_in ? 12'hb87 : _GEN_258; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_260 = 12'h104 == io_in ? 12'hfd7 : _GEN_259; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_261 = 12'h105 == io_in ? 12'hcc6 : _GEN_260; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_262 = 12'h106 == io_in ? 12'h8bb : _GEN_261; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_263 = 12'h107 == io_in ? 12'hced : _GEN_262; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_264 = 12'h108 == io_in ? 12'hb58 : _GEN_263; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_265 = 12'h109 == io_in ? 12'h278 : _GEN_264; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_266 = 12'h10a == io_in ? 12'hce6 : _GEN_265; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_267 = 12'h10b == io_in ? 12'h5d6 : _GEN_266; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_268 = 12'h10c == io_in ? 12'h3d : _GEN_267; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_269 = 12'h10d == io_in ? 12'h8e4 : _GEN_268; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_270 = 12'h10e == io_in ? 12'h81a : _GEN_269; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_271 = 12'h10f == io_in ? 12'h1b4 : _GEN_270; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_272 = 12'h110 == io_in ? 12'hf1a : _GEN_271; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_273 = 12'h111 == io_in ? 12'hbb : _GEN_272; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_274 = 12'h112 == io_in ? 12'h746 : _GEN_273; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_275 = 12'h113 == io_in ? 12'h529 : _GEN_274; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_276 = 12'h114 == io_in ? 12'hde7 : _GEN_275; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_277 = 12'h115 == io_in ? 12'hc9b : _GEN_276; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_278 = 12'h116 == io_in ? 12'h7aa : _GEN_277; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_279 = 12'h117 == io_in ? 12'h7d : _GEN_278; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_280 = 12'h118 == io_in ? 12'hb19 : _GEN_279; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_281 = 12'h119 == io_in ? 12'hed4 : _GEN_280; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_282 = 12'h11a == io_in ? 12'hd60 : _GEN_281; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_283 = 12'h11b == io_in ? 12'hbce : _GEN_282; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_284 = 12'h11c == io_in ? 12'h8f7 : _GEN_283; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_285 = 12'h11d == io_in ? 12'h374 : _GEN_284; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_286 = 12'h11e == io_in ? 12'h24d : _GEN_285; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_287 = 12'h11f == io_in ? 12'h44a : _GEN_286; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_288 = 12'h120 == io_in ? 12'hf9f : _GEN_287; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_289 = 12'h121 == io_in ? 12'h2a : _GEN_288; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_290 = 12'h122 == io_in ? 12'hacb : _GEN_289; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_291 = 12'h123 == io_in ? 12'h124 : _GEN_290; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_292 = 12'h124 == io_in ? 12'h74e : _GEN_291; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_293 = 12'h125 == io_in ? 12'h4a2 : _GEN_292; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_294 = 12'h126 == io_in ? 12'hd6f : _GEN_293; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_295 = 12'h127 == io_in ? 12'h18e : _GEN_294; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_296 = 12'h128 == io_in ? 12'h298 : _GEN_295; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_297 = 12'h129 == io_in ? 12'h63c : _GEN_296; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_298 = 12'h12a == io_in ? 12'h4f8 : _GEN_297; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_299 = 12'h12b == io_in ? 12'hbef : _GEN_298; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_300 = 12'h12c == io_in ? 12'hb17 : _GEN_299; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_301 = 12'h12d == io_in ? 12'hede : _GEN_300; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_302 = 12'h12e == io_in ? 12'hb12 : _GEN_301; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_303 = 12'h12f == io_in ? 12'hb42 : _GEN_302; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_304 = 12'h130 == io_in ? 12'hfe1 : _GEN_303; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_305 = 12'h131 == io_in ? 12'h6ce : _GEN_304; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_306 = 12'h132 == io_in ? 12'h2d4 : _GEN_305; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_307 = 12'h133 == io_in ? 12'h24 : _GEN_306; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_308 = 12'h134 == io_in ? 12'h62 : _GEN_307; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_309 = 12'h135 == io_in ? 12'ha8c : _GEN_308; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_310 = 12'h136 == io_in ? 12'h644 : _GEN_309; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_311 = 12'h137 == io_in ? 12'h4f4 : _GEN_310; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_312 = 12'h138 == io_in ? 12'h78b : _GEN_311; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_313 = 12'h139 == io_in ? 12'h75d : _GEN_312; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_314 = 12'h13a == io_in ? 12'h391 : _GEN_313; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_315 = 12'h13b == io_in ? 12'haa1 : _GEN_314; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_316 = 12'h13c == io_in ? 12'h9de : _GEN_315; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_317 = 12'h13d == io_in ? 12'h101 : _GEN_316; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_318 = 12'h13e == io_in ? 12'hef8 : _GEN_317; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_319 = 12'h13f == io_in ? 12'h1c : _GEN_318; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_320 = 12'h140 == io_in ? 12'he82 : _GEN_319; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_321 = 12'h141 == io_in ? 12'h1dd : _GEN_320; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_322 = 12'h142 == io_in ? 12'h513 : _GEN_321; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_323 = 12'h143 == io_in ? 12'h7fd : _GEN_322; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_324 = 12'h144 == io_in ? 12'ha36 : _GEN_323; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_325 = 12'h145 == io_in ? 12'h216 : _GEN_324; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_326 = 12'h146 == io_in ? 12'hf08 : _GEN_325; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_327 = 12'h147 == io_in ? 12'hdfc : _GEN_326; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_328 = 12'h148 == io_in ? 12'hed5 : _GEN_327; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_329 = 12'h149 == io_in ? 12'h352 : _GEN_328; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_330 = 12'h14a == io_in ? 12'h46b : _GEN_329; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_331 = 12'h14b == io_in ? 12'haf3 : _GEN_330; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_332 = 12'h14c == io_in ? 12'h790 : _GEN_331; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_333 = 12'h14d == io_in ? 12'h43a : _GEN_332; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_334 = 12'h14e == io_in ? 12'h502 : _GEN_333; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_335 = 12'h14f == io_in ? 12'h6cb : _GEN_334; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_336 = 12'h150 == io_in ? 12'hff9 : _GEN_335; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_337 = 12'h151 == io_in ? 12'h207 : _GEN_336; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_338 = 12'h152 == io_in ? 12'h312 : _GEN_337; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_339 = 12'h153 == io_in ? 12'h291 : _GEN_338; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_340 = 12'h154 == io_in ? 12'h10a : _GEN_339; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_341 = 12'h155 == io_in ? 12'h664 : _GEN_340; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_342 = 12'h156 == io_in ? 12'h310 : _GEN_341; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_343 = 12'h157 == io_in ? 12'hb02 : _GEN_342; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_344 = 12'h158 == io_in ? 12'hd19 : _GEN_343; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_345 = 12'h159 == io_in ? 12'h6c4 : _GEN_344; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_346 = 12'h15a == io_in ? 12'h265 : _GEN_345; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_347 = 12'h15b == io_in ? 12'hc5 : _GEN_346; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_348 = 12'h15c == io_in ? 12'h332 : _GEN_347; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_349 = 12'h15d == io_in ? 12'hf6c : _GEN_348; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_350 = 12'h15e == io_in ? 12'h6c : _GEN_349; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_351 = 12'h15f == io_in ? 12'h416 : _GEN_350; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_352 = 12'h160 == io_in ? 12'hfd0 : _GEN_351; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_353 = 12'h161 == io_in ? 12'h289 : _GEN_352; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_354 = 12'h162 == io_in ? 12'h448 : _GEN_353; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_355 = 12'h163 == io_in ? 12'h66c : _GEN_354; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_356 = 12'h164 == io_in ? 12'h7a9 : _GEN_355; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_357 = 12'h165 == io_in ? 12'h270 : _GEN_356; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_358 = 12'h166 == io_in ? 12'ha3f : _GEN_357; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_359 = 12'h167 == io_in ? 12'h6f7 : _GEN_358; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_360 = 12'h168 == io_in ? 12'h832 : _GEN_359; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_361 = 12'h169 == io_in ? 12'h8f9 : _GEN_360; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_362 = 12'h16a == io_in ? 12'h397 : _GEN_361; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_363 = 12'h16b == io_in ? 12'h37f : _GEN_362; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_364 = 12'h16c == io_in ? 12'h662 : _GEN_363; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_365 = 12'h16d == io_in ? 12'h516 : _GEN_364; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_366 = 12'h16e == io_in ? 12'he0d : _GEN_365; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_367 = 12'h16f == io_in ? 12'h430 : _GEN_366; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_368 = 12'h170 == io_in ? 12'h71 : _GEN_367; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_369 = 12'h171 == io_in ? 12'h6c3 : _GEN_368; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_370 = 12'h172 == io_in ? 12'h16e : _GEN_369; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_371 = 12'h173 == io_in ? 12'h7ab : _GEN_370; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_372 = 12'h174 == io_in ? 12'h311 : _GEN_371; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_373 = 12'h175 == io_in ? 12'h195 : _GEN_372; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_374 = 12'h176 == io_in ? 12'h334 : _GEN_373; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_375 = 12'h177 == io_in ? 12'h77a : _GEN_374; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_376 = 12'h178 == io_in ? 12'h1ea : _GEN_375; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_377 = 12'h179 == io_in ? 12'haf4 : _GEN_376; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_378 = 12'h17a == io_in ? 12'h518 : _GEN_377; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_379 = 12'h17b == io_in ? 12'h1ce : _GEN_378; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_380 = 12'h17c == io_in ? 12'h9e : _GEN_379; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_381 = 12'h17d == io_in ? 12'h49c : _GEN_380; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_382 = 12'h17e == io_in ? 12'h342 : _GEN_381; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_383 = 12'h17f == io_in ? 12'hb32 : _GEN_382; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_384 = 12'h180 == io_in ? 12'hbd0 : _GEN_383; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_385 = 12'h181 == io_in ? 12'ha59 : _GEN_384; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_386 = 12'h182 == io_in ? 12'h3e2 : _GEN_385; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_387 = 12'h183 == io_in ? 12'h3c1 : _GEN_386; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_388 = 12'h184 == io_in ? 12'hda9 : _GEN_387; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_389 = 12'h185 == io_in ? 12'h553 : _GEN_388; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_390 = 12'h186 == io_in ? 12'h95f : _GEN_389; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_391 = 12'h187 == io_in ? 12'h30a : _GEN_390; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_392 = 12'h188 == io_in ? 12'h82f : _GEN_391; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_393 = 12'h189 == io_in ? 12'h49c : _GEN_392; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_394 = 12'h18a == io_in ? 12'h3b8 : _GEN_393; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_395 = 12'h18b == io_in ? 12'hb03 : _GEN_394; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_396 = 12'h18c == io_in ? 12'h142 : _GEN_395; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_397 = 12'h18d == io_in ? 12'hcc6 : _GEN_396; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_398 = 12'h18e == io_in ? 12'h822 : _GEN_397; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_399 = 12'h18f == io_in ? 12'hcec : _GEN_398; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_400 = 12'h190 == io_in ? 12'hb4c : _GEN_399; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_401 = 12'h191 == io_in ? 12'h3f9 : _GEN_400; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_402 = 12'h192 == io_in ? 12'hff5 : _GEN_401; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_403 = 12'h193 == io_in ? 12'he94 : _GEN_402; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_404 = 12'h194 == io_in ? 12'hd60 : _GEN_403; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_405 = 12'h195 == io_in ? 12'h150 : _GEN_404; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_406 = 12'h196 == io_in ? 12'haca : _GEN_405; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_407 = 12'h197 == io_in ? 12'hee8 : _GEN_406; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_408 = 12'h198 == io_in ? 12'hb28 : _GEN_407; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_409 = 12'h199 == io_in ? 12'h21d : _GEN_408; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_410 = 12'h19a == io_in ? 12'h289 : _GEN_409; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_411 = 12'h19b == io_in ? 12'h6aa : _GEN_410; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_412 = 12'h19c == io_in ? 12'h595 : _GEN_411; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_413 = 12'h19d == io_in ? 12'h28b : _GEN_412; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_414 = 12'h19e == io_in ? 12'hacd : _GEN_413; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_415 = 12'h19f == io_in ? 12'hdb6 : _GEN_414; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_416 = 12'h1a0 == io_in ? 12'h101 : _GEN_415; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_417 = 12'h1a1 == io_in ? 12'hec4 : _GEN_416; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_418 = 12'h1a2 == io_in ? 12'h4e1 : _GEN_417; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_419 = 12'h1a3 == io_in ? 12'hba3 : _GEN_418; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_420 = 12'h1a4 == io_in ? 12'hbf8 : _GEN_419; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_421 = 12'h1a5 == io_in ? 12'h2b1 : _GEN_420; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_422 = 12'h1a6 == io_in ? 12'h564 : _GEN_421; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_423 = 12'h1a7 == io_in ? 12'h830 : _GEN_422; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_424 = 12'h1a8 == io_in ? 12'hd6d : _GEN_423; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_425 = 12'h1a9 == io_in ? 12'h76c : _GEN_424; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_426 = 12'h1aa == io_in ? 12'h3ff : _GEN_425; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_427 = 12'h1ab == io_in ? 12'h6d6 : _GEN_426; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_428 = 12'h1ac == io_in ? 12'h42d : _GEN_427; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_429 = 12'h1ad == io_in ? 12'h335 : _GEN_428; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_430 = 12'h1ae == io_in ? 12'hdad : _GEN_429; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_431 = 12'h1af == io_in ? 12'h1bf : _GEN_430; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_432 = 12'h1b0 == io_in ? 12'hf8 : _GEN_431; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_433 = 12'h1b1 == io_in ? 12'h280 : _GEN_432; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_434 = 12'h1b2 == io_in ? 12'h143 : _GEN_433; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_435 = 12'h1b3 == io_in ? 12'h1ae : _GEN_434; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_436 = 12'h1b4 == io_in ? 12'h4dd : _GEN_435; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_437 = 12'h1b5 == io_in ? 12'hbcd : _GEN_436; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_438 = 12'h1b6 == io_in ? 12'h7a9 : _GEN_437; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_439 = 12'h1b7 == io_in ? 12'hfc3 : _GEN_438; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_440 = 12'h1b8 == io_in ? 12'h6b1 : _GEN_439; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_441 = 12'h1b9 == io_in ? 12'h41e : _GEN_440; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_442 = 12'h1ba == io_in ? 12'he78 : _GEN_441; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_443 = 12'h1bb == io_in ? 12'h5c6 : _GEN_442; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_444 = 12'h1bc == io_in ? 12'h305 : _GEN_443; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_445 = 12'h1bd == io_in ? 12'hcf0 : _GEN_444; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_446 = 12'h1be == io_in ? 12'h66e : _GEN_445; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_447 = 12'h1bf == io_in ? 12'h46d : _GEN_446; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_448 = 12'h1c0 == io_in ? 12'hc71 : _GEN_447; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_449 = 12'h1c1 == io_in ? 12'h694 : _GEN_448; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_450 = 12'h1c2 == io_in ? 12'hee4 : _GEN_449; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_451 = 12'h1c3 == io_in ? 12'hb71 : _GEN_450; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_452 = 12'h1c4 == io_in ? 12'hfc5 : _GEN_451; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_453 = 12'h1c5 == io_in ? 12'h159 : _GEN_452; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_454 = 12'h1c6 == io_in ? 12'h464 : _GEN_453; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_455 = 12'h1c7 == io_in ? 12'h48c : _GEN_454; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_456 = 12'h1c8 == io_in ? 12'h542 : _GEN_455; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_457 = 12'h1c9 == io_in ? 12'h58f : _GEN_456; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_458 = 12'h1ca == io_in ? 12'h8fc : _GEN_457; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_459 = 12'h1cb == io_in ? 12'h367 : _GEN_458; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_460 = 12'h1cc == io_in ? 12'h985 : _GEN_459; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_461 = 12'h1cd == io_in ? 12'hcd2 : _GEN_460; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_462 = 12'h1ce == io_in ? 12'h78e : _GEN_461; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_463 = 12'h1cf == io_in ? 12'h56b : _GEN_462; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_464 = 12'h1d0 == io_in ? 12'h594 : _GEN_463; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_465 = 12'h1d1 == io_in ? 12'hfdd : _GEN_464; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_466 = 12'h1d2 == io_in ? 12'hcae : _GEN_465; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_467 = 12'h1d3 == io_in ? 12'hc12 : _GEN_466; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_468 = 12'h1d4 == io_in ? 12'h37c : _GEN_467; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_469 = 12'h1d5 == io_in ? 12'ha18 : _GEN_468; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_470 = 12'h1d6 == io_in ? 12'hd72 : _GEN_469; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_471 = 12'h1d7 == io_in ? 12'hbaf : _GEN_470; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_472 = 12'h1d8 == io_in ? 12'he8c : _GEN_471; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_473 = 12'h1d9 == io_in ? 12'h975 : _GEN_472; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_474 = 12'h1da == io_in ? 12'h10f : _GEN_473; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_475 = 12'h1db == io_in ? 12'hb43 : _GEN_474; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_476 = 12'h1dc == io_in ? 12'h3de : _GEN_475; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_477 = 12'h1dd == io_in ? 12'h573 : _GEN_476; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_478 = 12'h1de == io_in ? 12'h23a : _GEN_477; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_479 = 12'h1df == io_in ? 12'hce4 : _GEN_478; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_480 = 12'h1e0 == io_in ? 12'h5f3 : _GEN_479; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_481 = 12'h1e1 == io_in ? 12'hd80 : _GEN_480; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_482 = 12'h1e2 == io_in ? 12'h182 : _GEN_481; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_483 = 12'h1e3 == io_in ? 12'h1bc : _GEN_482; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_484 = 12'h1e4 == io_in ? 12'h20 : _GEN_483; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_485 = 12'h1e5 == io_in ? 12'h612 : _GEN_484; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_486 = 12'h1e6 == io_in ? 12'hd44 : _GEN_485; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_487 = 12'h1e7 == io_in ? 12'ha36 : _GEN_486; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_488 = 12'h1e8 == io_in ? 12'h319 : _GEN_487; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_489 = 12'h1e9 == io_in ? 12'h6e0 : _GEN_488; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_490 = 12'h1ea == io_in ? 12'he4d : _GEN_489; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_491 = 12'h1eb == io_in ? 12'hf76 : _GEN_490; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_492 = 12'h1ec == io_in ? 12'hfc : _GEN_491; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_493 = 12'h1ed == io_in ? 12'h512 : _GEN_492; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_494 = 12'h1ee == io_in ? 12'h26c : _GEN_493; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_495 = 12'h1ef == io_in ? 12'hc82 : _GEN_494; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_496 = 12'h1f0 == io_in ? 12'h606 : _GEN_495; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_497 = 12'h1f1 == io_in ? 12'hca7 : _GEN_496; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_498 = 12'h1f2 == io_in ? 12'h6db : _GEN_497; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_499 = 12'h1f3 == io_in ? 12'h50b : _GEN_498; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_500 = 12'h1f4 == io_in ? 12'h41d : _GEN_499; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_501 = 12'h1f5 == io_in ? 12'h67c : _GEN_500; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_502 = 12'h1f6 == io_in ? 12'haf4 : _GEN_501; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_503 = 12'h1f7 == io_in ? 12'h7cc : _GEN_502; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_504 = 12'h1f8 == io_in ? 12'he35 : _GEN_503; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_505 = 12'h1f9 == io_in ? 12'h7cb : _GEN_504; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_506 = 12'h1fa == io_in ? 12'hcc1 : _GEN_505; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_507 = 12'h1fb == io_in ? 12'h932 : _GEN_506; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_508 = 12'h1fc == io_in ? 12'h865 : _GEN_507; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_509 = 12'h1fd == io_in ? 12'h678 : _GEN_508; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_510 = 12'h1fe == io_in ? 12'haf2 : _GEN_509; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_511 = 12'h1ff == io_in ? 12'h6c8 : _GEN_510; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_512 = 12'h200 == io_in ? 12'h81b : _GEN_511; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_513 = 12'h201 == io_in ? 12'hf5c : _GEN_512; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_514 = 12'h202 == io_in ? 12'hdfd : _GEN_513; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_515 = 12'h203 == io_in ? 12'h7cc : _GEN_514; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_516 = 12'h204 == io_in ? 12'h343 : _GEN_515; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_517 = 12'h205 == io_in ? 12'h347 : _GEN_516; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_518 = 12'h206 == io_in ? 12'h8c8 : _GEN_517; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_519 = 12'h207 == io_in ? 12'h611 : _GEN_518; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_520 = 12'h208 == io_in ? 12'hda7 : _GEN_519; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_521 = 12'h209 == io_in ? 12'h13c : _GEN_520; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_522 = 12'h20a == io_in ? 12'haa3 : _GEN_521; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_523 = 12'h20b == io_in ? 12'h35f : _GEN_522; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_524 = 12'h20c == io_in ? 12'h954 : _GEN_523; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_525 = 12'h20d == io_in ? 12'hb80 : _GEN_524; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_526 = 12'h20e == io_in ? 12'hb52 : _GEN_525; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_527 = 12'h20f == io_in ? 12'ha44 : _GEN_526; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_528 = 12'h210 == io_in ? 12'hce3 : _GEN_527; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_529 = 12'h211 == io_in ? 12'h679 : _GEN_528; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_530 = 12'h212 == io_in ? 12'h68b : _GEN_529; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_531 = 12'h213 == io_in ? 12'h9a4 : _GEN_530; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_532 = 12'h214 == io_in ? 12'hb3b : _GEN_531; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_533 = 12'h215 == io_in ? 12'hf75 : _GEN_532; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_534 = 12'h216 == io_in ? 12'hdd : _GEN_533; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_535 = 12'h217 == io_in ? 12'hc1b : _GEN_534; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_536 = 12'h218 == io_in ? 12'h1b9 : _GEN_535; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_537 = 12'h219 == io_in ? 12'hc0a : _GEN_536; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_538 = 12'h21a == io_in ? 12'ha72 : _GEN_537; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_539 = 12'h21b == io_in ? 12'h7f0 : _GEN_538; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_540 = 12'h21c == io_in ? 12'h85b : _GEN_539; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_541 = 12'h21d == io_in ? 12'h47a : _GEN_540; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_542 = 12'h21e == io_in ? 12'hd43 : _GEN_541; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_543 = 12'h21f == io_in ? 12'h246 : _GEN_542; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_544 = 12'h220 == io_in ? 12'hc0c : _GEN_543; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_545 = 12'h221 == io_in ? 12'h2cc : _GEN_544; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_546 = 12'h222 == io_in ? 12'h143 : _GEN_545; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_547 = 12'h223 == io_in ? 12'hd37 : _GEN_546; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_548 = 12'h224 == io_in ? 12'h4af : _GEN_547; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_549 = 12'h225 == io_in ? 12'h143 : _GEN_548; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_550 = 12'h226 == io_in ? 12'h7e8 : _GEN_549; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_551 = 12'h227 == io_in ? 12'h9b5 : _GEN_550; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_552 = 12'h228 == io_in ? 12'h9ed : _GEN_551; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_553 = 12'h229 == io_in ? 12'h45f : _GEN_552; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_554 = 12'h22a == io_in ? 12'he15 : _GEN_553; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_555 = 12'h22b == io_in ? 12'hc76 : _GEN_554; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_556 = 12'h22c == io_in ? 12'h4e8 : _GEN_555; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_557 = 12'h22d == io_in ? 12'hb5d : _GEN_556; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_558 = 12'h22e == io_in ? 12'hb99 : _GEN_557; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_559 = 12'h22f == io_in ? 12'h28a : _GEN_558; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_560 = 12'h230 == io_in ? 12'hf22 : _GEN_559; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_561 = 12'h231 == io_in ? 12'h574 : _GEN_560; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_562 = 12'h232 == io_in ? 12'hdc8 : _GEN_561; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_563 = 12'h233 == io_in ? 12'hc4a : _GEN_562; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_564 = 12'h234 == io_in ? 12'h474 : _GEN_563; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_565 = 12'h235 == io_in ? 12'h731 : _GEN_564; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_566 = 12'h236 == io_in ? 12'h1bb : _GEN_565; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_567 = 12'h237 == io_in ? 12'h9eb : _GEN_566; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_568 = 12'h238 == io_in ? 12'h6a2 : _GEN_567; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_569 = 12'h239 == io_in ? 12'h9fc : _GEN_568; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_570 = 12'h23a == io_in ? 12'h3f4 : _GEN_569; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_571 = 12'h23b == io_in ? 12'he84 : _GEN_570; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_572 = 12'h23c == io_in ? 12'h3ee : _GEN_571; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_573 = 12'h23d == io_in ? 12'hdec : _GEN_572; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_574 = 12'h23e == io_in ? 12'h864 : _GEN_573; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_575 = 12'h23f == io_in ? 12'h783 : _GEN_574; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_576 = 12'h240 == io_in ? 12'h116 : _GEN_575; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_577 = 12'h241 == io_in ? 12'hb92 : _GEN_576; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_578 = 12'h242 == io_in ? 12'h638 : _GEN_577; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_579 = 12'h243 == io_in ? 12'hd8c : _GEN_578; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_580 = 12'h244 == io_in ? 12'h40f : _GEN_579; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_581 = 12'h245 == io_in ? 12'h6fe : _GEN_580; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_582 = 12'h246 == io_in ? 12'h77c : _GEN_581; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_583 = 12'h247 == io_in ? 12'h6a : _GEN_582; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_584 = 12'h248 == io_in ? 12'hc09 : _GEN_583; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_585 = 12'h249 == io_in ? 12'hf53 : _GEN_584; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_586 = 12'h24a == io_in ? 12'h2c3 : _GEN_585; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_587 = 12'h24b == io_in ? 12'h472 : _GEN_586; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_588 = 12'h24c == io_in ? 12'h10b : _GEN_587; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_589 = 12'h24d == io_in ? 12'h5ce : _GEN_588; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_590 = 12'h24e == io_in ? 12'hc2a : _GEN_589; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_591 = 12'h24f == io_in ? 12'h8c3 : _GEN_590; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_592 = 12'h250 == io_in ? 12'h8aa : _GEN_591; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_593 = 12'h251 == io_in ? 12'h551 : _GEN_592; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_594 = 12'h252 == io_in ? 12'hf5d : _GEN_593; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_595 = 12'h253 == io_in ? 12'h279 : _GEN_594; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_596 = 12'h254 == io_in ? 12'hcd1 : _GEN_595; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_597 = 12'h255 == io_in ? 12'h7a7 : _GEN_596; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_598 = 12'h256 == io_in ? 12'h34d : _GEN_597; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_599 = 12'h257 == io_in ? 12'h15b : _GEN_598; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_600 = 12'h258 == io_in ? 12'h6ac : _GEN_599; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_601 = 12'h259 == io_in ? 12'h98a : _GEN_600; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_602 = 12'h25a == io_in ? 12'h4d6 : _GEN_601; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_603 = 12'h25b == io_in ? 12'hb12 : _GEN_602; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_604 = 12'h25c == io_in ? 12'hb7f : _GEN_603; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_605 = 12'h25d == io_in ? 12'h1b7 : _GEN_604; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_606 = 12'h25e == io_in ? 12'hbf3 : _GEN_605; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_607 = 12'h25f == io_in ? 12'hf1d : _GEN_606; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_608 = 12'h260 == io_in ? 12'h827 : _GEN_607; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_609 = 12'h261 == io_in ? 12'hc66 : _GEN_608; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_610 = 12'h262 == io_in ? 12'h85c : _GEN_609; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_611 = 12'h263 == io_in ? 12'h805 : _GEN_610; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_612 = 12'h264 == io_in ? 12'h4f4 : _GEN_611; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_613 = 12'h265 == io_in ? 12'hb78 : _GEN_612; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_614 = 12'h266 == io_in ? 12'h935 : _GEN_613; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_615 = 12'h267 == io_in ? 12'h72c : _GEN_614; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_616 = 12'h268 == io_in ? 12'h5db : _GEN_615; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_617 = 12'h269 == io_in ? 12'h770 : _GEN_616; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_618 = 12'h26a == io_in ? 12'h7ce : _GEN_617; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_619 = 12'h26b == io_in ? 12'hce5 : _GEN_618; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_620 = 12'h26c == io_in ? 12'h834 : _GEN_619; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_621 = 12'h26d == io_in ? 12'h6a2 : _GEN_620; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_622 = 12'h26e == io_in ? 12'h809 : _GEN_621; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_623 = 12'h26f == io_in ? 12'h404 : _GEN_622; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_624 = 12'h270 == io_in ? 12'h9f : _GEN_623; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_625 = 12'h271 == io_in ? 12'h204 : _GEN_624; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_626 = 12'h272 == io_in ? 12'h89a : _GEN_625; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_627 = 12'h273 == io_in ? 12'h87d : _GEN_626; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_628 = 12'h274 == io_in ? 12'h1ed : _GEN_627; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_629 = 12'h275 == io_in ? 12'h33d : _GEN_628; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_630 = 12'h276 == io_in ? 12'h927 : _GEN_629; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_631 = 12'h277 == io_in ? 12'hdee : _GEN_630; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_632 = 12'h278 == io_in ? 12'h456 : _GEN_631; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_633 = 12'h279 == io_in ? 12'h97d : _GEN_632; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_634 = 12'h27a == io_in ? 12'h978 : _GEN_633; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_635 = 12'h27b == io_in ? 12'h35f : _GEN_634; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_636 = 12'h27c == io_in ? 12'h63a : _GEN_635; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_637 = 12'h27d == io_in ? 12'h441 : _GEN_636; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_638 = 12'h27e == io_in ? 12'h932 : _GEN_637; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_639 = 12'h27f == io_in ? 12'h3c5 : _GEN_638; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_640 = 12'h280 == io_in ? 12'hb09 : _GEN_639; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_641 = 12'h281 == io_in ? 12'h64 : _GEN_640; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_642 = 12'h282 == io_in ? 12'heb8 : _GEN_641; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_643 = 12'h283 == io_in ? 12'h152 : _GEN_642; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_644 = 12'h284 == io_in ? 12'h75d : _GEN_643; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_645 = 12'h285 == io_in ? 12'h7a7 : _GEN_644; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_646 = 12'h286 == io_in ? 12'h9e6 : _GEN_645; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_647 = 12'h287 == io_in ? 12'hfcb : _GEN_646; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_648 = 12'h288 == io_in ? 12'hb76 : _GEN_647; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_649 = 12'h289 == io_in ? 12'h8e7 : _GEN_648; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_650 = 12'h28a == io_in ? 12'he96 : _GEN_649; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_651 = 12'h28b == io_in ? 12'h6cc : _GEN_650; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_652 = 12'h28c == io_in ? 12'h6fa : _GEN_651; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_653 = 12'h28d == io_in ? 12'hb9b : _GEN_652; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_654 = 12'h28e == io_in ? 12'h635 : _GEN_653; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_655 = 12'h28f == io_in ? 12'h21 : _GEN_654; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_656 = 12'h290 == io_in ? 12'hd92 : _GEN_655; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_657 = 12'h291 == io_in ? 12'hfed : _GEN_656; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_658 = 12'h292 == io_in ? 12'h76f : _GEN_657; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_659 = 12'h293 == io_in ? 12'h33f : _GEN_658; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_660 = 12'h294 == io_in ? 12'hde1 : _GEN_659; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_661 = 12'h295 == io_in ? 12'h9f6 : _GEN_660; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_662 = 12'h296 == io_in ? 12'ha3 : _GEN_661; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_663 = 12'h297 == io_in ? 12'h22a : _GEN_662; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_664 = 12'h298 == io_in ? 12'h138 : _GEN_663; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_665 = 12'h299 == io_in ? 12'hfd7 : _GEN_664; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_666 = 12'h29a == io_in ? 12'h47f : _GEN_665; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_667 = 12'h29b == io_in ? 12'h566 : _GEN_666; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_668 = 12'h29c == io_in ? 12'hf75 : _GEN_667; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_669 = 12'h29d == io_in ? 12'hb02 : _GEN_668; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_670 = 12'h29e == io_in ? 12'hf86 : _GEN_669; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_671 = 12'h29f == io_in ? 12'h4e0 : _GEN_670; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_672 = 12'h2a0 == io_in ? 12'h76e : _GEN_671; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_673 = 12'h2a1 == io_in ? 12'h402 : _GEN_672; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_674 = 12'h2a2 == io_in ? 12'h71d : _GEN_673; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_675 = 12'h2a3 == io_in ? 12'h76f : _GEN_674; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_676 = 12'h2a4 == io_in ? 12'h111 : _GEN_675; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_677 = 12'h2a5 == io_in ? 12'hf1 : _GEN_676; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_678 = 12'h2a6 == io_in ? 12'hd1f : _GEN_677; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_679 = 12'h2a7 == io_in ? 12'h70f : _GEN_678; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_680 = 12'h2a8 == io_in ? 12'h563 : _GEN_679; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_681 = 12'h2a9 == io_in ? 12'h8e1 : _GEN_680; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_682 = 12'h2aa == io_in ? 12'h24f : _GEN_681; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_683 = 12'h2ab == io_in ? 12'he29 : _GEN_682; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_684 = 12'h2ac == io_in ? 12'hbe1 : _GEN_683; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_685 = 12'h2ad == io_in ? 12'h653 : _GEN_684; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_686 = 12'h2ae == io_in ? 12'h2d2 : _GEN_685; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_687 = 12'h2af == io_in ? 12'h3e0 : _GEN_686; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_688 = 12'h2b0 == io_in ? 12'h172 : _GEN_687; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_689 = 12'h2b1 == io_in ? 12'h79a : _GEN_688; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_690 = 12'h2b2 == io_in ? 12'h4d2 : _GEN_689; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_691 = 12'h2b3 == io_in ? 12'h826 : _GEN_690; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_692 = 12'h2b4 == io_in ? 12'h809 : _GEN_691; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_693 = 12'h2b5 == io_in ? 12'hb3e : _GEN_692; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_694 = 12'h2b6 == io_in ? 12'h621 : _GEN_693; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_695 = 12'h2b7 == io_in ? 12'ha48 : _GEN_694; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_696 = 12'h2b8 == io_in ? 12'h631 : _GEN_695; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_697 = 12'h2b9 == io_in ? 12'hfb5 : _GEN_696; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_698 = 12'h2ba == io_in ? 12'h28a : _GEN_697; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_699 = 12'h2bb == io_in ? 12'hff9 : _GEN_698; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_700 = 12'h2bc == io_in ? 12'h2e9 : _GEN_699; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_701 = 12'h2bd == io_in ? 12'h6b1 : _GEN_700; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_702 = 12'h2be == io_in ? 12'hc52 : _GEN_701; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_703 = 12'h2bf == io_in ? 12'h241 : _GEN_702; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_704 = 12'h2c0 == io_in ? 12'h5d2 : _GEN_703; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_705 = 12'h2c1 == io_in ? 12'h59a : _GEN_704; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_706 = 12'h2c2 == io_in ? 12'h9b3 : _GEN_705; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_707 = 12'h2c3 == io_in ? 12'hf89 : _GEN_706; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_708 = 12'h2c4 == io_in ? 12'hfc2 : _GEN_707; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_709 = 12'h2c5 == io_in ? 12'h438 : _GEN_708; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_710 = 12'h2c6 == io_in ? 12'h614 : _GEN_709; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_711 = 12'h2c7 == io_in ? 12'h5f3 : _GEN_710; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_712 = 12'h2c8 == io_in ? 12'h8b5 : _GEN_711; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_713 = 12'h2c9 == io_in ? 12'h12f : _GEN_712; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_714 = 12'h2ca == io_in ? 12'h1e9 : _GEN_713; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_715 = 12'h2cb == io_in ? 12'h1ab : _GEN_714; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_716 = 12'h2cc == io_in ? 12'h9f6 : _GEN_715; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_717 = 12'h2cd == io_in ? 12'haa : _GEN_716; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_718 = 12'h2ce == io_in ? 12'hfa8 : _GEN_717; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_719 = 12'h2cf == io_in ? 12'h430 : _GEN_718; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_720 = 12'h2d0 == io_in ? 12'h552 : _GEN_719; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_721 = 12'h2d1 == io_in ? 12'hd1a : _GEN_720; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_722 = 12'h2d2 == io_in ? 12'hb77 : _GEN_721; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_723 = 12'h2d3 == io_in ? 12'h305 : _GEN_722; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_724 = 12'h2d4 == io_in ? 12'h290 : _GEN_723; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_725 = 12'h2d5 == io_in ? 12'hc38 : _GEN_724; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_726 = 12'h2d6 == io_in ? 12'hb98 : _GEN_725; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_727 = 12'h2d7 == io_in ? 12'hdf6 : _GEN_726; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_728 = 12'h2d8 == io_in ? 12'h55f : _GEN_727; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_729 = 12'h2d9 == io_in ? 12'hcc9 : _GEN_728; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_730 = 12'h2da == io_in ? 12'h442 : _GEN_729; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_731 = 12'h2db == io_in ? 12'hb75 : _GEN_730; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_732 = 12'h2dc == io_in ? 12'hfb4 : _GEN_731; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_733 = 12'h2dd == io_in ? 12'h3f7 : _GEN_732; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_734 = 12'h2de == io_in ? 12'h61a : _GEN_733; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_735 = 12'h2df == io_in ? 12'h8e8 : _GEN_734; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_736 = 12'h2e0 == io_in ? 12'h428 : _GEN_735; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_737 = 12'h2e1 == io_in ? 12'h589 : _GEN_736; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_738 = 12'h2e2 == io_in ? 12'hcdb : _GEN_737; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_739 = 12'h2e3 == io_in ? 12'h5f8 : _GEN_738; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_740 = 12'h2e4 == io_in ? 12'hc0e : _GEN_739; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_741 = 12'h2e5 == io_in ? 12'h979 : _GEN_740; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_742 = 12'h2e6 == io_in ? 12'h5da : _GEN_741; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_743 = 12'h2e7 == io_in ? 12'h5ed : _GEN_742; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_744 = 12'h2e8 == io_in ? 12'hce7 : _GEN_743; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_745 = 12'h2e9 == io_in ? 12'hd86 : _GEN_744; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_746 = 12'h2ea == io_in ? 12'h43c : _GEN_745; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_747 = 12'h2eb == io_in ? 12'he6a : _GEN_746; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_748 = 12'h2ec == io_in ? 12'h63f : _GEN_747; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_749 = 12'h2ed == io_in ? 12'hbc7 : _GEN_748; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_750 = 12'h2ee == io_in ? 12'h3f5 : _GEN_749; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_751 = 12'h2ef == io_in ? 12'hc78 : _GEN_750; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_752 = 12'h2f0 == io_in ? 12'hd03 : _GEN_751; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_753 = 12'h2f1 == io_in ? 12'hadf : _GEN_752; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_754 = 12'h2f2 == io_in ? 12'h2d7 : _GEN_753; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_755 = 12'h2f3 == io_in ? 12'h21a : _GEN_754; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_756 = 12'h2f4 == io_in ? 12'hcd5 : _GEN_755; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_757 = 12'h2f5 == io_in ? 12'haa2 : _GEN_756; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_758 = 12'h2f6 == io_in ? 12'h87c : _GEN_757; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_759 = 12'h2f7 == io_in ? 12'h92a : _GEN_758; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_760 = 12'h2f8 == io_in ? 12'hdeb : _GEN_759; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_761 = 12'h2f9 == io_in ? 12'h460 : _GEN_760; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_762 = 12'h2fa == io_in ? 12'h6b3 : _GEN_761; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_763 = 12'h2fb == io_in ? 12'ha82 : _GEN_762; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_764 = 12'h2fc == io_in ? 12'ha30 : _GEN_763; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_765 = 12'h2fd == io_in ? 12'habd : _GEN_764; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_766 = 12'h2fe == io_in ? 12'haf8 : _GEN_765; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_767 = 12'h2ff == io_in ? 12'h8dc : _GEN_766; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_768 = 12'h300 == io_in ? 12'hc59 : _GEN_767; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_769 = 12'h301 == io_in ? 12'hdd3 : _GEN_768; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_770 = 12'h302 == io_in ? 12'h15f : _GEN_769; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_771 = 12'h303 == io_in ? 12'h845 : _GEN_770; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_772 = 12'h304 == io_in ? 12'h540 : _GEN_771; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_773 = 12'h305 == io_in ? 12'h7f6 : _GEN_772; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_774 = 12'h306 == io_in ? 12'h6ee : _GEN_773; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_775 = 12'h307 == io_in ? 12'h4a : _GEN_774; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_776 = 12'h308 == io_in ? 12'h796 : _GEN_775; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_777 = 12'h309 == io_in ? 12'h24f : _GEN_776; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_778 = 12'h30a == io_in ? 12'he93 : _GEN_777; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_779 = 12'h30b == io_in ? 12'h7b8 : _GEN_778; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_780 = 12'h30c == io_in ? 12'h7f2 : _GEN_779; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_781 = 12'h30d == io_in ? 12'h1a7 : _GEN_780; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_782 = 12'h30e == io_in ? 12'h383 : _GEN_781; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_783 = 12'h30f == io_in ? 12'h3f8 : _GEN_782; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_784 = 12'h310 == io_in ? 12'ha7a : _GEN_783; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_785 = 12'h311 == io_in ? 12'h831 : _GEN_784; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_786 = 12'h312 == io_in ? 12'h68a : _GEN_785; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_787 = 12'h313 == io_in ? 12'h1e : _GEN_786; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_788 = 12'h314 == io_in ? 12'h298 : _GEN_787; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_789 = 12'h315 == io_in ? 12'h451 : _GEN_788; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_790 = 12'h316 == io_in ? 12'haec : _GEN_789; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_791 = 12'h317 == io_in ? 12'h401 : _GEN_790; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_792 = 12'h318 == io_in ? 12'h9a3 : _GEN_791; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_793 = 12'h319 == io_in ? 12'h3f5 : _GEN_792; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_794 = 12'h31a == io_in ? 12'h1fa : _GEN_793; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_795 = 12'h31b == io_in ? 12'haec : _GEN_794; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_796 = 12'h31c == io_in ? 12'h495 : _GEN_795; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_797 = 12'h31d == io_in ? 12'h3fd : _GEN_796; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_798 = 12'h31e == io_in ? 12'ha65 : _GEN_797; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_799 = 12'h31f == io_in ? 12'hc0d : _GEN_798; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_800 = 12'h320 == io_in ? 12'he92 : _GEN_799; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_801 = 12'h321 == io_in ? 12'h961 : _GEN_800; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_802 = 12'h322 == io_in ? 12'heec : _GEN_801; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_803 = 12'h323 == io_in ? 12'h140 : _GEN_802; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_804 = 12'h324 == io_in ? 12'hdee : _GEN_803; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_805 = 12'h325 == io_in ? 12'h2f1 : _GEN_804; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_806 = 12'h326 == io_in ? 12'he10 : _GEN_805; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_807 = 12'h327 == io_in ? 12'h94 : _GEN_806; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_808 = 12'h328 == io_in ? 12'h5fe : _GEN_807; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_809 = 12'h329 == io_in ? 12'h502 : _GEN_808; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_810 = 12'h32a == io_in ? 12'h57b : _GEN_809; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_811 = 12'h32b == io_in ? 12'h2f3 : _GEN_810; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_812 = 12'h32c == io_in ? 12'h386 : _GEN_811; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_813 = 12'h32d == io_in ? 12'h13e : _GEN_812; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_814 = 12'h32e == io_in ? 12'h51c : _GEN_813; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_815 = 12'h32f == io_in ? 12'h82f : _GEN_814; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_816 = 12'h330 == io_in ? 12'h905 : _GEN_815; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_817 = 12'h331 == io_in ? 12'h32c : _GEN_816; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_818 = 12'h332 == io_in ? 12'h1eb : _GEN_817; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_819 = 12'h333 == io_in ? 12'h464 : _GEN_818; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_820 = 12'h334 == io_in ? 12'hffe : _GEN_819; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_821 = 12'h335 == io_in ? 12'hb29 : _GEN_820; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_822 = 12'h336 == io_in ? 12'h233 : _GEN_821; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_823 = 12'h337 == io_in ? 12'h1b0 : _GEN_822; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_824 = 12'h338 == io_in ? 12'hc66 : _GEN_823; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_825 = 12'h339 == io_in ? 12'h55a : _GEN_824; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_826 = 12'h33a == io_in ? 12'h63f : _GEN_825; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_827 = 12'h33b == io_in ? 12'he82 : _GEN_826; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_828 = 12'h33c == io_in ? 12'h66e : _GEN_827; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_829 = 12'h33d == io_in ? 12'he32 : _GEN_828; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_830 = 12'h33e == io_in ? 12'h24a : _GEN_829; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_831 = 12'h33f == io_in ? 12'h64c : _GEN_830; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_832 = 12'h340 == io_in ? 12'h763 : _GEN_831; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_833 = 12'h341 == io_in ? 12'h2cb : _GEN_832; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_834 = 12'h342 == io_in ? 12'h8e9 : _GEN_833; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_835 = 12'h343 == io_in ? 12'hf2b : _GEN_834; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_836 = 12'h344 == io_in ? 12'h160 : _GEN_835; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_837 = 12'h345 == io_in ? 12'h6fb : _GEN_836; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_838 = 12'h346 == io_in ? 12'h86e : _GEN_837; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_839 = 12'h347 == io_in ? 12'h20d : _GEN_838; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_840 = 12'h348 == io_in ? 12'hc4f : _GEN_839; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_841 = 12'h349 == io_in ? 12'he17 : _GEN_840; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_842 = 12'h34a == io_in ? 12'hfe9 : _GEN_841; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_843 = 12'h34b == io_in ? 12'hf75 : _GEN_842; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_844 = 12'h34c == io_in ? 12'h88e : _GEN_843; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_845 = 12'h34d == io_in ? 12'hd29 : _GEN_844; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_846 = 12'h34e == io_in ? 12'h43 : _GEN_845; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_847 = 12'h34f == io_in ? 12'h45f : _GEN_846; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_848 = 12'h350 == io_in ? 12'h851 : _GEN_847; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_849 = 12'h351 == io_in ? 12'h659 : _GEN_848; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_850 = 12'h352 == io_in ? 12'h812 : _GEN_849; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_851 = 12'h353 == io_in ? 12'h108 : _GEN_850; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_852 = 12'h354 == io_in ? 12'h25f : _GEN_851; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_853 = 12'h355 == io_in ? 12'hdbc : _GEN_852; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_854 = 12'h356 == io_in ? 12'ha9c : _GEN_853; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_855 = 12'h357 == io_in ? 12'he87 : _GEN_854; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_856 = 12'h358 == io_in ? 12'hd5d : _GEN_855; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_857 = 12'h359 == io_in ? 12'h86c : _GEN_856; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_858 = 12'h35a == io_in ? 12'heff : _GEN_857; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_859 = 12'h35b == io_in ? 12'h40a : _GEN_858; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_860 = 12'h35c == io_in ? 12'hae2 : _GEN_859; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_861 = 12'h35d == io_in ? 12'h848 : _GEN_860; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_862 = 12'h35e == io_in ? 12'h76a : _GEN_861; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_863 = 12'h35f == io_in ? 12'h64e : _GEN_862; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_864 = 12'h360 == io_in ? 12'h9ae : _GEN_863; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_865 = 12'h361 == io_in ? 12'h2b0 : _GEN_864; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_866 = 12'h362 == io_in ? 12'h393 : _GEN_865; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_867 = 12'h363 == io_in ? 12'hbeb : _GEN_866; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_868 = 12'h364 == io_in ? 12'h9c5 : _GEN_867; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_869 = 12'h365 == io_in ? 12'hfcc : _GEN_868; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_870 = 12'h366 == io_in ? 12'hf18 : _GEN_869; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_871 = 12'h367 == io_in ? 12'h35 : _GEN_870; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_872 = 12'h368 == io_in ? 12'h2cc : _GEN_871; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_873 = 12'h369 == io_in ? 12'hc84 : _GEN_872; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_874 = 12'h36a == io_in ? 12'h4ac : _GEN_873; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_875 = 12'h36b == io_in ? 12'h292 : _GEN_874; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_876 = 12'h36c == io_in ? 12'ha67 : _GEN_875; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_877 = 12'h36d == io_in ? 12'h4e9 : _GEN_876; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_878 = 12'h36e == io_in ? 12'ha47 : _GEN_877; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_879 = 12'h36f == io_in ? 12'he16 : _GEN_878; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_880 = 12'h370 == io_in ? 12'hf45 : _GEN_879; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_881 = 12'h371 == io_in ? 12'h1c9 : _GEN_880; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_882 = 12'h372 == io_in ? 12'h1b : _GEN_881; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_883 = 12'h373 == io_in ? 12'h72d : _GEN_882; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_884 = 12'h374 == io_in ? 12'hde6 : _GEN_883; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_885 = 12'h375 == io_in ? 12'hc68 : _GEN_884; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_886 = 12'h376 == io_in ? 12'h294 : _GEN_885; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_887 = 12'h377 == io_in ? 12'h501 : _GEN_886; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_888 = 12'h378 == io_in ? 12'h205 : _GEN_887; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_889 = 12'h379 == io_in ? 12'h25d : _GEN_888; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_890 = 12'h37a == io_in ? 12'h4ac : _GEN_889; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_891 = 12'h37b == io_in ? 12'h844 : _GEN_890; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_892 = 12'h37c == io_in ? 12'hdc3 : _GEN_891; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_893 = 12'h37d == io_in ? 12'hb2b : _GEN_892; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_894 = 12'h37e == io_in ? 12'h114 : _GEN_893; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_895 = 12'h37f == io_in ? 12'hfc2 : _GEN_894; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_896 = 12'h380 == io_in ? 12'h465 : _GEN_895; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_897 = 12'h381 == io_in ? 12'h5a2 : _GEN_896; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_898 = 12'h382 == io_in ? 12'h16b : _GEN_897; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_899 = 12'h383 == io_in ? 12'hf56 : _GEN_898; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_900 = 12'h384 == io_in ? 12'hf42 : _GEN_899; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_901 = 12'h385 == io_in ? 12'heb6 : _GEN_900; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_902 = 12'h386 == io_in ? 12'h7d1 : _GEN_901; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_903 = 12'h387 == io_in ? 12'h269 : _GEN_902; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_904 = 12'h388 == io_in ? 12'h8c4 : _GEN_903; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_905 = 12'h389 == io_in ? 12'h2c9 : _GEN_904; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_906 = 12'h38a == io_in ? 12'ha31 : _GEN_905; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_907 = 12'h38b == io_in ? 12'hf9c : _GEN_906; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_908 = 12'h38c == io_in ? 12'hbb1 : _GEN_907; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_909 = 12'h38d == io_in ? 12'hb8 : _GEN_908; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_910 = 12'h38e == io_in ? 12'ha9a : _GEN_909; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_911 = 12'h38f == io_in ? 12'hecc : _GEN_910; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_912 = 12'h390 == io_in ? 12'hea3 : _GEN_911; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_913 = 12'h391 == io_in ? 12'hfcc : _GEN_912; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_914 = 12'h392 == io_in ? 12'hdbf : _GEN_913; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_915 = 12'h393 == io_in ? 12'h94d : _GEN_914; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_916 = 12'h394 == io_in ? 12'h6 : _GEN_915; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_917 = 12'h395 == io_in ? 12'h30e : _GEN_916; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_918 = 12'h396 == io_in ? 12'h118 : _GEN_917; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_919 = 12'h397 == io_in ? 12'h1e3 : _GEN_918; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_920 = 12'h398 == io_in ? 12'h30d : _GEN_919; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_921 = 12'h399 == io_in ? 12'ha86 : _GEN_920; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_922 = 12'h39a == io_in ? 12'h494 : _GEN_921; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_923 = 12'h39b == io_in ? 12'h6fd : _GEN_922; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_924 = 12'h39c == io_in ? 12'hf73 : _GEN_923; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_925 = 12'h39d == io_in ? 12'h9db : _GEN_924; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_926 = 12'h39e == io_in ? 12'h2b : _GEN_925; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_927 = 12'h39f == io_in ? 12'h674 : _GEN_926; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_928 = 12'h3a0 == io_in ? 12'hc1b : _GEN_927; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_929 = 12'h3a1 == io_in ? 12'h19f : _GEN_928; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_930 = 12'h3a2 == io_in ? 12'hf9 : _GEN_929; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_931 = 12'h3a3 == io_in ? 12'h383 : _GEN_930; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_932 = 12'h3a4 == io_in ? 12'h7c6 : _GEN_931; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_933 = 12'h3a5 == io_in ? 12'h999 : _GEN_932; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_934 = 12'h3a6 == io_in ? 12'hb24 : _GEN_933; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_935 = 12'h3a7 == io_in ? 12'ha86 : _GEN_934; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_936 = 12'h3a8 == io_in ? 12'h550 : _GEN_935; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_937 = 12'h3a9 == io_in ? 12'h592 : _GEN_936; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_938 = 12'h3aa == io_in ? 12'h98 : _GEN_937; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_939 = 12'h3ab == io_in ? 12'h404 : _GEN_938; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_940 = 12'h3ac == io_in ? 12'h49f : _GEN_939; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_941 = 12'h3ad == io_in ? 12'h7e9 : _GEN_940; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_942 = 12'h3ae == io_in ? 12'he84 : _GEN_941; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_943 = 12'h3af == io_in ? 12'h292 : _GEN_942; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_944 = 12'h3b0 == io_in ? 12'hb84 : _GEN_943; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_945 = 12'h3b1 == io_in ? 12'hd32 : _GEN_944; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_946 = 12'h3b2 == io_in ? 12'he3a : _GEN_945; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_947 = 12'h3b3 == io_in ? 12'h39a : _GEN_946; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_948 = 12'h3b4 == io_in ? 12'h6b6 : _GEN_947; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_949 = 12'h3b5 == io_in ? 12'hf53 : _GEN_948; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_950 = 12'h3b6 == io_in ? 12'h57a : _GEN_949; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_951 = 12'h3b7 == io_in ? 12'hf73 : _GEN_950; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_952 = 12'h3b8 == io_in ? 12'h2fd : _GEN_951; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_953 = 12'h3b9 == io_in ? 12'hccc : _GEN_952; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_954 = 12'h3ba == io_in ? 12'h721 : _GEN_953; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_955 = 12'h3bb == io_in ? 12'h435 : _GEN_954; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_956 = 12'h3bc == io_in ? 12'h79d : _GEN_955; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_957 = 12'h3bd == io_in ? 12'h17 : _GEN_956; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_958 = 12'h3be == io_in ? 12'h97a : _GEN_957; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_959 = 12'h3bf == io_in ? 12'h288 : _GEN_958; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_960 = 12'h3c0 == io_in ? 12'h5e : _GEN_959; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_961 = 12'h3c1 == io_in ? 12'h31c : _GEN_960; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_962 = 12'h3c2 == io_in ? 12'h2db : _GEN_961; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_963 = 12'h3c3 == io_in ? 12'h337 : _GEN_962; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_964 = 12'h3c4 == io_in ? 12'hfb6 : _GEN_963; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_965 = 12'h3c5 == io_in ? 12'ha76 : _GEN_964; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_966 = 12'h3c6 == io_in ? 12'h7cf : _GEN_965; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_967 = 12'h3c7 == io_in ? 12'hea6 : _GEN_966; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_968 = 12'h3c8 == io_in ? 12'hde6 : _GEN_967; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_969 = 12'h3c9 == io_in ? 12'h3e0 : _GEN_968; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_970 = 12'h3ca == io_in ? 12'he17 : _GEN_969; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_971 = 12'h3cb == io_in ? 12'hf82 : _GEN_970; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_972 = 12'h3cc == io_in ? 12'hc15 : _GEN_971; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_973 = 12'h3cd == io_in ? 12'h9d2 : _GEN_972; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_974 = 12'h3ce == io_in ? 12'h41f : _GEN_973; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_975 = 12'h3cf == io_in ? 12'h3cc : _GEN_974; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_976 = 12'h3d0 == io_in ? 12'h998 : _GEN_975; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_977 = 12'h3d1 == io_in ? 12'hd1b : _GEN_976; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_978 = 12'h3d2 == io_in ? 12'h180 : _GEN_977; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_979 = 12'h3d3 == io_in ? 12'h26a : _GEN_978; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_980 = 12'h3d4 == io_in ? 12'h483 : _GEN_979; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_981 = 12'h3d5 == io_in ? 12'hb77 : _GEN_980; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_982 = 12'h3d6 == io_in ? 12'h872 : _GEN_981; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_983 = 12'h3d7 == io_in ? 12'hfb0 : _GEN_982; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_984 = 12'h3d8 == io_in ? 12'heb2 : _GEN_983; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_985 = 12'h3d9 == io_in ? 12'h99e : _GEN_984; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_986 = 12'h3da == io_in ? 12'hc60 : _GEN_985; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_987 = 12'h3db == io_in ? 12'h54b : _GEN_986; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_988 = 12'h3dc == io_in ? 12'heb6 : _GEN_987; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_989 = 12'h3dd == io_in ? 12'h793 : _GEN_988; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_990 = 12'h3de == io_in ? 12'hb5b : _GEN_989; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_991 = 12'h3df == io_in ? 12'h5b6 : _GEN_990; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_992 = 12'h3e0 == io_in ? 12'h4e9 : _GEN_991; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_993 = 12'h3e1 == io_in ? 12'h99f : _GEN_992; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_994 = 12'h3e2 == io_in ? 12'h21 : _GEN_993; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_995 = 12'h3e3 == io_in ? 12'ha5a : _GEN_994; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_996 = 12'h3e4 == io_in ? 12'h35f : _GEN_995; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_997 = 12'h3e5 == io_in ? 12'h785 : _GEN_996; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_998 = 12'h3e6 == io_in ? 12'hb7a : _GEN_997; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_999 = 12'h3e7 == io_in ? 12'h5e8 : _GEN_998; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1000 = 12'h3e8 == io_in ? 12'habd : _GEN_999; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1001 = 12'h3e9 == io_in ? 12'hca : _GEN_1000; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1002 = 12'h3ea == io_in ? 12'h5aa : _GEN_1001; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1003 = 12'h3eb == io_in ? 12'h53 : _GEN_1002; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1004 = 12'h3ec == io_in ? 12'hb8f : _GEN_1003; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1005 = 12'h3ed == io_in ? 12'h156 : _GEN_1004; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1006 = 12'h3ee == io_in ? 12'h4a2 : _GEN_1005; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1007 = 12'h3ef == io_in ? 12'hc01 : _GEN_1006; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1008 = 12'h3f0 == io_in ? 12'hd44 : _GEN_1007; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1009 = 12'h3f1 == io_in ? 12'h5c : _GEN_1008; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1010 = 12'h3f2 == io_in ? 12'h7cc : _GEN_1009; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1011 = 12'h3f3 == io_in ? 12'heb6 : _GEN_1010; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1012 = 12'h3f4 == io_in ? 12'h973 : _GEN_1011; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1013 = 12'h3f5 == io_in ? 12'h5b8 : _GEN_1012; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1014 = 12'h3f6 == io_in ? 12'h680 : _GEN_1013; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1015 = 12'h3f7 == io_in ? 12'hdae : _GEN_1014; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1016 = 12'h3f8 == io_in ? 12'hfaa : _GEN_1015; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1017 = 12'h3f9 == io_in ? 12'hb71 : _GEN_1016; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1018 = 12'h3fa == io_in ? 12'h6e1 : _GEN_1017; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1019 = 12'h3fb == io_in ? 12'h24a : _GEN_1018; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1020 = 12'h3fc == io_in ? 12'h654 : _GEN_1019; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1021 = 12'h3fd == io_in ? 12'hbbe : _GEN_1020; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1022 = 12'h3fe == io_in ? 12'h6ae : _GEN_1021; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1023 = 12'h3ff == io_in ? 12'h9aa : _GEN_1022; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1024 = 12'h400 == io_in ? 12'h6a3 : _GEN_1023; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1025 = 12'h401 == io_in ? 12'hbe7 : _GEN_1024; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1026 = 12'h402 == io_in ? 12'h903 : _GEN_1025; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1027 = 12'h403 == io_in ? 12'h7d : _GEN_1026; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1028 = 12'h404 == io_in ? 12'h149 : _GEN_1027; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1029 = 12'h405 == io_in ? 12'hbe7 : _GEN_1028; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1030 = 12'h406 == io_in ? 12'h8c7 : _GEN_1029; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1031 = 12'h407 == io_in ? 12'h49 : _GEN_1030; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1032 = 12'h408 == io_in ? 12'hff : _GEN_1031; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1033 = 12'h409 == io_in ? 12'h6cd : _GEN_1032; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1034 = 12'h40a == io_in ? 12'h1e : _GEN_1033; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1035 = 12'h40b == io_in ? 12'hb7f : _GEN_1034; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1036 = 12'h40c == io_in ? 12'h5e3 : _GEN_1035; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1037 = 12'h40d == io_in ? 12'haec : _GEN_1036; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1038 = 12'h40e == io_in ? 12'h604 : _GEN_1037; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1039 = 12'h40f == io_in ? 12'h1b4 : _GEN_1038; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1040 = 12'h410 == io_in ? 12'hd85 : _GEN_1039; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1041 = 12'h411 == io_in ? 12'h870 : _GEN_1040; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1042 = 12'h412 == io_in ? 12'hb71 : _GEN_1041; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1043 = 12'h413 == io_in ? 12'h8ae : _GEN_1042; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1044 = 12'h414 == io_in ? 12'h8b1 : _GEN_1043; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1045 = 12'h415 == io_in ? 12'hc47 : _GEN_1044; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1046 = 12'h416 == io_in ? 12'hb99 : _GEN_1045; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1047 = 12'h417 == io_in ? 12'hdef : _GEN_1046; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1048 = 12'h418 == io_in ? 12'h81b : _GEN_1047; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1049 = 12'h419 == io_in ? 12'h9dd : _GEN_1048; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1050 = 12'h41a == io_in ? 12'hce0 : _GEN_1049; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1051 = 12'h41b == io_in ? 12'h733 : _GEN_1050; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1052 = 12'h41c == io_in ? 12'h850 : _GEN_1051; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1053 = 12'h41d == io_in ? 12'h422 : _GEN_1052; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1054 = 12'h41e == io_in ? 12'h319 : _GEN_1053; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1055 = 12'h41f == io_in ? 12'hf5e : _GEN_1054; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1056 = 12'h420 == io_in ? 12'h46a : _GEN_1055; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1057 = 12'h421 == io_in ? 12'hbab : _GEN_1056; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1058 = 12'h422 == io_in ? 12'h3da : _GEN_1057; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1059 = 12'h423 == io_in ? 12'h573 : _GEN_1058; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1060 = 12'h424 == io_in ? 12'hd47 : _GEN_1059; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1061 = 12'h425 == io_in ? 12'h8dd : _GEN_1060; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1062 = 12'h426 == io_in ? 12'h2a5 : _GEN_1061; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1063 = 12'h427 == io_in ? 12'h18c : _GEN_1062; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1064 = 12'h428 == io_in ? 12'hacc : _GEN_1063; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1065 = 12'h429 == io_in ? 12'hca6 : _GEN_1064; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1066 = 12'h42a == io_in ? 12'hf5e : _GEN_1065; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1067 = 12'h42b == io_in ? 12'h93b : _GEN_1066; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1068 = 12'h42c == io_in ? 12'h8cb : _GEN_1067; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1069 = 12'h42d == io_in ? 12'h544 : _GEN_1068; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1070 = 12'h42e == io_in ? 12'hbe3 : _GEN_1069; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1071 = 12'h42f == io_in ? 12'hb58 : _GEN_1070; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1072 = 12'h430 == io_in ? 12'hda4 : _GEN_1071; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1073 = 12'h431 == io_in ? 12'hdfa : _GEN_1072; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1074 = 12'h432 == io_in ? 12'hf04 : _GEN_1073; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1075 = 12'h433 == io_in ? 12'h852 : _GEN_1074; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1076 = 12'h434 == io_in ? 12'h311 : _GEN_1075; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1077 = 12'h435 == io_in ? 12'h5cc : _GEN_1076; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1078 = 12'h436 == io_in ? 12'h831 : _GEN_1077; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1079 = 12'h437 == io_in ? 12'h5d5 : _GEN_1078; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1080 = 12'h438 == io_in ? 12'he3 : _GEN_1079; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1081 = 12'h439 == io_in ? 12'h241 : _GEN_1080; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1082 = 12'h43a == io_in ? 12'h7c1 : _GEN_1081; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1083 = 12'h43b == io_in ? 12'hd66 : _GEN_1082; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1084 = 12'h43c == io_in ? 12'h4ba : _GEN_1083; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1085 = 12'h43d == io_in ? 12'hd42 : _GEN_1084; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1086 = 12'h43e == io_in ? 12'h6a4 : _GEN_1085; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1087 = 12'h43f == io_in ? 12'h798 : _GEN_1086; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1088 = 12'h440 == io_in ? 12'h3b8 : _GEN_1087; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1089 = 12'h441 == io_in ? 12'hdf : _GEN_1088; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1090 = 12'h442 == io_in ? 12'h475 : _GEN_1089; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1091 = 12'h443 == io_in ? 12'h7f7 : _GEN_1090; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1092 = 12'h444 == io_in ? 12'hc62 : _GEN_1091; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1093 = 12'h445 == io_in ? 12'h799 : _GEN_1092; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1094 = 12'h446 == io_in ? 12'h4fc : _GEN_1093; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1095 = 12'h447 == io_in ? 12'h736 : _GEN_1094; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1096 = 12'h448 == io_in ? 12'h50c : _GEN_1095; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1097 = 12'h449 == io_in ? 12'h3c2 : _GEN_1096; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1098 = 12'h44a == io_in ? 12'h41a : _GEN_1097; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1099 = 12'h44b == io_in ? 12'hd4e : _GEN_1098; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1100 = 12'h44c == io_in ? 12'h142 : _GEN_1099; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1101 = 12'h44d == io_in ? 12'h476 : _GEN_1100; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1102 = 12'h44e == io_in ? 12'hfc8 : _GEN_1101; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1103 = 12'h44f == io_in ? 12'hf46 : _GEN_1102; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1104 = 12'h450 == io_in ? 12'h6c1 : _GEN_1103; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1105 = 12'h451 == io_in ? 12'h2d6 : _GEN_1104; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1106 = 12'h452 == io_in ? 12'h7d3 : _GEN_1105; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1107 = 12'h453 == io_in ? 12'hc25 : _GEN_1106; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1108 = 12'h454 == io_in ? 12'he62 : _GEN_1107; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1109 = 12'h455 == io_in ? 12'he76 : _GEN_1108; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1110 = 12'h456 == io_in ? 12'h786 : _GEN_1109; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1111 = 12'h457 == io_in ? 12'h229 : _GEN_1110; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1112 = 12'h458 == io_in ? 12'h13d : _GEN_1111; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1113 = 12'h459 == io_in ? 12'hdfa : _GEN_1112; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1114 = 12'h45a == io_in ? 12'h9dc : _GEN_1113; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1115 = 12'h45b == io_in ? 12'h511 : _GEN_1114; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1116 = 12'h45c == io_in ? 12'h6a4 : _GEN_1115; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1117 = 12'h45d == io_in ? 12'h819 : _GEN_1116; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1118 = 12'h45e == io_in ? 12'h89c : _GEN_1117; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1119 = 12'h45f == io_in ? 12'hc6a : _GEN_1118; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1120 = 12'h460 == io_in ? 12'h909 : _GEN_1119; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1121 = 12'h461 == io_in ? 12'h491 : _GEN_1120; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1122 = 12'h462 == io_in ? 12'h3b4 : _GEN_1121; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1123 = 12'h463 == io_in ? 12'he63 : _GEN_1122; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1124 = 12'h464 == io_in ? 12'h193 : _GEN_1123; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1125 = 12'h465 == io_in ? 12'h396 : _GEN_1124; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1126 = 12'h466 == io_in ? 12'h2a9 : _GEN_1125; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1127 = 12'h467 == io_in ? 12'h194 : _GEN_1126; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1128 = 12'h468 == io_in ? 12'hb11 : _GEN_1127; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1129 = 12'h469 == io_in ? 12'h83e : _GEN_1128; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1130 = 12'h46a == io_in ? 12'hdb8 : _GEN_1129; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1131 = 12'h46b == io_in ? 12'h390 : _GEN_1130; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1132 = 12'h46c == io_in ? 12'hab2 : _GEN_1131; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1133 = 12'h46d == io_in ? 12'hfc3 : _GEN_1132; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1134 = 12'h46e == io_in ? 12'h8b2 : _GEN_1133; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1135 = 12'h46f == io_in ? 12'h8cf : _GEN_1134; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1136 = 12'h470 == io_in ? 12'h92b : _GEN_1135; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1137 = 12'h471 == io_in ? 12'h7bd : _GEN_1136; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1138 = 12'h472 == io_in ? 12'hcaf : _GEN_1137; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1139 = 12'h473 == io_in ? 12'hdeb : _GEN_1138; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1140 = 12'h474 == io_in ? 12'h18b : _GEN_1139; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1141 = 12'h475 == io_in ? 12'h1a8 : _GEN_1140; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1142 = 12'h476 == io_in ? 12'hf43 : _GEN_1141; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1143 = 12'h477 == io_in ? 12'h4a4 : _GEN_1142; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1144 = 12'h478 == io_in ? 12'h850 : _GEN_1143; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1145 = 12'h479 == io_in ? 12'he27 : _GEN_1144; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1146 = 12'h47a == io_in ? 12'h299 : _GEN_1145; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1147 = 12'h47b == io_in ? 12'h6b8 : _GEN_1146; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1148 = 12'h47c == io_in ? 12'h7af : _GEN_1147; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1149 = 12'h47d == io_in ? 12'h822 : _GEN_1148; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1150 = 12'h47e == io_in ? 12'h7c7 : _GEN_1149; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1151 = 12'h47f == io_in ? 12'h3c9 : _GEN_1150; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1152 = 12'h480 == io_in ? 12'hc22 : _GEN_1151; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1153 = 12'h481 == io_in ? 12'h351 : _GEN_1152; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1154 = 12'h482 == io_in ? 12'hf7c : _GEN_1153; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1155 = 12'h483 == io_in ? 12'h977 : _GEN_1154; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1156 = 12'h484 == io_in ? 12'h34c : _GEN_1155; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1157 = 12'h485 == io_in ? 12'h586 : _GEN_1156; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1158 = 12'h486 == io_in ? 12'hc4 : _GEN_1157; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1159 = 12'h487 == io_in ? 12'h7d6 : _GEN_1158; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1160 = 12'h488 == io_in ? 12'h80b : _GEN_1159; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1161 = 12'h489 == io_in ? 12'ha72 : _GEN_1160; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1162 = 12'h48a == io_in ? 12'hc9d : _GEN_1161; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1163 = 12'h48b == io_in ? 12'h873 : _GEN_1162; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1164 = 12'h48c == io_in ? 12'hed : _GEN_1163; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1165 = 12'h48d == io_in ? 12'h1e4 : _GEN_1164; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1166 = 12'h48e == io_in ? 12'h9f1 : _GEN_1165; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1167 = 12'h48f == io_in ? 12'ha55 : _GEN_1166; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1168 = 12'h490 == io_in ? 12'hd7e : _GEN_1167; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1169 = 12'h491 == io_in ? 12'hd78 : _GEN_1168; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1170 = 12'h492 == io_in ? 12'hff : _GEN_1169; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1171 = 12'h493 == io_in ? 12'h576 : _GEN_1170; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1172 = 12'h494 == io_in ? 12'hd7b : _GEN_1171; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1173 = 12'h495 == io_in ? 12'h823 : _GEN_1172; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1174 = 12'h496 == io_in ? 12'h74 : _GEN_1173; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1175 = 12'h497 == io_in ? 12'h97 : _GEN_1174; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1176 = 12'h498 == io_in ? 12'h86 : _GEN_1175; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1177 = 12'h499 == io_in ? 12'h501 : _GEN_1176; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1178 = 12'h49a == io_in ? 12'h8da : _GEN_1177; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1179 = 12'h49b == io_in ? 12'h4c3 : _GEN_1178; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1180 = 12'h49c == io_in ? 12'ha73 : _GEN_1179; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1181 = 12'h49d == io_in ? 12'h7ec : _GEN_1180; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1182 = 12'h49e == io_in ? 12'hbec : _GEN_1181; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1183 = 12'h49f == io_in ? 12'h333 : _GEN_1182; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1184 = 12'h4a0 == io_in ? 12'h1a : _GEN_1183; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1185 = 12'h4a1 == io_in ? 12'hf2f : _GEN_1184; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1186 = 12'h4a2 == io_in ? 12'haf4 : _GEN_1185; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1187 = 12'h4a3 == io_in ? 12'h933 : _GEN_1186; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1188 = 12'h4a4 == io_in ? 12'h1cd : _GEN_1187; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1189 = 12'h4a5 == io_in ? 12'h6ce : _GEN_1188; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1190 = 12'h4a6 == io_in ? 12'h73c : _GEN_1189; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1191 = 12'h4a7 == io_in ? 12'hf38 : _GEN_1190; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1192 = 12'h4a8 == io_in ? 12'h64c : _GEN_1191; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1193 = 12'h4a9 == io_in ? 12'ha12 : _GEN_1192; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1194 = 12'h4aa == io_in ? 12'heb8 : _GEN_1193; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1195 = 12'h4ab == io_in ? 12'h5a0 : _GEN_1194; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1196 = 12'h4ac == io_in ? 12'hcff : _GEN_1195; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1197 = 12'h4ad == io_in ? 12'h3e8 : _GEN_1196; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1198 = 12'h4ae == io_in ? 12'h157 : _GEN_1197; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1199 = 12'h4af == io_in ? 12'h47e : _GEN_1198; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1200 = 12'h4b0 == io_in ? 12'hda4 : _GEN_1199; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1201 = 12'h4b1 == io_in ? 12'h99e : _GEN_1200; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1202 = 12'h4b2 == io_in ? 12'h42c : _GEN_1201; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1203 = 12'h4b3 == io_in ? 12'h18b : _GEN_1202; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1204 = 12'h4b4 == io_in ? 12'haf0 : _GEN_1203; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1205 = 12'h4b5 == io_in ? 12'h2d2 : _GEN_1204; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1206 = 12'h4b6 == io_in ? 12'h1c5 : _GEN_1205; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1207 = 12'h4b7 == io_in ? 12'he97 : _GEN_1206; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1208 = 12'h4b8 == io_in ? 12'h4ba : _GEN_1207; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1209 = 12'h4b9 == io_in ? 12'h4c0 : _GEN_1208; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1210 = 12'h4ba == io_in ? 12'h3b8 : _GEN_1209; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1211 = 12'h4bb == io_in ? 12'h526 : _GEN_1210; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1212 = 12'h4bc == io_in ? 12'h3b5 : _GEN_1211; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1213 = 12'h4bd == io_in ? 12'hc45 : _GEN_1212; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1214 = 12'h4be == io_in ? 12'haa9 : _GEN_1213; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1215 = 12'h4bf == io_in ? 12'hc61 : _GEN_1214; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1216 = 12'h4c0 == io_in ? 12'h73d : _GEN_1215; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1217 = 12'h4c1 == io_in ? 12'h940 : _GEN_1216; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1218 = 12'h4c2 == io_in ? 12'h713 : _GEN_1217; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1219 = 12'h4c3 == io_in ? 12'hbb9 : _GEN_1218; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1220 = 12'h4c4 == io_in ? 12'h652 : _GEN_1219; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1221 = 12'h4c5 == io_in ? 12'h591 : _GEN_1220; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1222 = 12'h4c6 == io_in ? 12'hebe : _GEN_1221; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1223 = 12'h4c7 == io_in ? 12'hd3a : _GEN_1222; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1224 = 12'h4c8 == io_in ? 12'h455 : _GEN_1223; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1225 = 12'h4c9 == io_in ? 12'had8 : _GEN_1224; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1226 = 12'h4ca == io_in ? 12'he6f : _GEN_1225; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1227 = 12'h4cb == io_in ? 12'haa0 : _GEN_1226; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1228 = 12'h4cc == io_in ? 12'h4c6 : _GEN_1227; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1229 = 12'h4cd == io_in ? 12'haaa : _GEN_1228; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1230 = 12'h4ce == io_in ? 12'hcb6 : _GEN_1229; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1231 = 12'h4cf == io_in ? 12'ha6a : _GEN_1230; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1232 = 12'h4d0 == io_in ? 12'hd94 : _GEN_1231; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1233 = 12'h4d1 == io_in ? 12'h6ea : _GEN_1232; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1234 = 12'h4d2 == io_in ? 12'hd58 : _GEN_1233; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1235 = 12'h4d3 == io_in ? 12'heca : _GEN_1234; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1236 = 12'h4d4 == io_in ? 12'h500 : _GEN_1235; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1237 = 12'h4d5 == io_in ? 12'ha1a : _GEN_1236; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1238 = 12'h4d6 == io_in ? 12'hb14 : _GEN_1237; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1239 = 12'h4d7 == io_in ? 12'hf43 : _GEN_1238; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1240 = 12'h4d8 == io_in ? 12'hf31 : _GEN_1239; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1241 = 12'h4d9 == io_in ? 12'hc12 : _GEN_1240; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1242 = 12'h4da == io_in ? 12'h990 : _GEN_1241; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1243 = 12'h4db == io_in ? 12'hb0e : _GEN_1242; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1244 = 12'h4dc == io_in ? 12'ha67 : _GEN_1243; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1245 = 12'h4dd == io_in ? 12'hdf3 : _GEN_1244; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1246 = 12'h4de == io_in ? 12'h795 : _GEN_1245; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1247 = 12'h4df == io_in ? 12'hb10 : _GEN_1246; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1248 = 12'h4e0 == io_in ? 12'hab5 : _GEN_1247; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1249 = 12'h4e1 == io_in ? 12'habd : _GEN_1248; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1250 = 12'h4e2 == io_in ? 12'hb86 : _GEN_1249; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1251 = 12'h4e3 == io_in ? 12'he49 : _GEN_1250; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1252 = 12'h4e4 == io_in ? 12'h305 : _GEN_1251; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1253 = 12'h4e5 == io_in ? 12'h150 : _GEN_1252; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1254 = 12'h4e6 == io_in ? 12'h3f2 : _GEN_1253; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1255 = 12'h4e7 == io_in ? 12'hcec : _GEN_1254; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1256 = 12'h4e8 == io_in ? 12'h7c1 : _GEN_1255; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1257 = 12'h4e9 == io_in ? 12'hac6 : _GEN_1256; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1258 = 12'h4ea == io_in ? 12'hbcc : _GEN_1257; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1259 = 12'h4eb == io_in ? 12'h999 : _GEN_1258; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1260 = 12'h4ec == io_in ? 12'h560 : _GEN_1259; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1261 = 12'h4ed == io_in ? 12'hecc : _GEN_1260; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1262 = 12'h4ee == io_in ? 12'heab : _GEN_1261; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1263 = 12'h4ef == io_in ? 12'hb06 : _GEN_1262; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1264 = 12'h4f0 == io_in ? 12'hbed : _GEN_1263; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1265 = 12'h4f1 == io_in ? 12'h91c : _GEN_1264; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1266 = 12'h4f2 == io_in ? 12'hb62 : _GEN_1265; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1267 = 12'h4f3 == io_in ? 12'h4b3 : _GEN_1266; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1268 = 12'h4f4 == io_in ? 12'h87e : _GEN_1267; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1269 = 12'h4f5 == io_in ? 12'h9be : _GEN_1268; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1270 = 12'h4f6 == io_in ? 12'ha54 : _GEN_1269; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1271 = 12'h4f7 == io_in ? 12'h50e : _GEN_1270; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1272 = 12'h4f8 == io_in ? 12'ha63 : _GEN_1271; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1273 = 12'h4f9 == io_in ? 12'h822 : _GEN_1272; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1274 = 12'h4fa == io_in ? 12'hd5c : _GEN_1273; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1275 = 12'h4fb == io_in ? 12'h8ab : _GEN_1274; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1276 = 12'h4fc == io_in ? 12'h684 : _GEN_1275; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1277 = 12'h4fd == io_in ? 12'h1f7 : _GEN_1276; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1278 = 12'h4fe == io_in ? 12'h7bb : _GEN_1277; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1279 = 12'h4ff == io_in ? 12'hbd4 : _GEN_1278; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1280 = 12'h500 == io_in ? 12'he0e : _GEN_1279; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1281 = 12'h501 == io_in ? 12'h5a9 : _GEN_1280; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1282 = 12'h502 == io_in ? 12'h7d8 : _GEN_1281; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1283 = 12'h503 == io_in ? 12'h844 : _GEN_1282; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1284 = 12'h504 == io_in ? 12'hbce : _GEN_1283; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1285 = 12'h505 == io_in ? 12'h810 : _GEN_1284; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1286 = 12'h506 == io_in ? 12'h802 : _GEN_1285; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1287 = 12'h507 == io_in ? 12'hf42 : _GEN_1286; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1288 = 12'h508 == io_in ? 12'h5ef : _GEN_1287; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1289 = 12'h509 == io_in ? 12'h1f5 : _GEN_1288; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1290 = 12'h50a == io_in ? 12'h804 : _GEN_1289; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1291 = 12'h50b == io_in ? 12'h17 : _GEN_1290; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1292 = 12'h50c == io_in ? 12'h6a : _GEN_1291; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1293 = 12'h50d == io_in ? 12'h748 : _GEN_1292; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1294 = 12'h50e == io_in ? 12'habd : _GEN_1293; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1295 = 12'h50f == io_in ? 12'h765 : _GEN_1294; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1296 = 12'h510 == io_in ? 12'h25c : _GEN_1295; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1297 = 12'h511 == io_in ? 12'hc6a : _GEN_1296; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1298 = 12'h512 == io_in ? 12'h143 : _GEN_1297; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1299 = 12'h513 == io_in ? 12'haf : _GEN_1298; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1300 = 12'h514 == io_in ? 12'h2b : _GEN_1299; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1301 = 12'h515 == io_in ? 12'h157 : _GEN_1300; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1302 = 12'h516 == io_in ? 12'h9be : _GEN_1301; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1303 = 12'h517 == io_in ? 12'hd2a : _GEN_1302; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1304 = 12'h518 == io_in ? 12'hb9a : _GEN_1303; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1305 = 12'h519 == io_in ? 12'h42b : _GEN_1304; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1306 = 12'h51a == io_in ? 12'h25f : _GEN_1305; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1307 = 12'h51b == io_in ? 12'hfe : _GEN_1306; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1308 = 12'h51c == io_in ? 12'h6ac : _GEN_1307; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1309 = 12'h51d == io_in ? 12'h86e : _GEN_1308; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1310 = 12'h51e == io_in ? 12'h5a : _GEN_1309; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1311 = 12'h51f == io_in ? 12'h3fc : _GEN_1310; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1312 = 12'h520 == io_in ? 12'h682 : _GEN_1311; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1313 = 12'h521 == io_in ? 12'h50f : _GEN_1312; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1314 = 12'h522 == io_in ? 12'h4f6 : _GEN_1313; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1315 = 12'h523 == io_in ? 12'h848 : _GEN_1314; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1316 = 12'h524 == io_in ? 12'hfe6 : _GEN_1315; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1317 = 12'h525 == io_in ? 12'hc1b : _GEN_1316; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1318 = 12'h526 == io_in ? 12'h676 : _GEN_1317; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1319 = 12'h527 == io_in ? 12'he82 : _GEN_1318; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1320 = 12'h528 == io_in ? 12'ha8a : _GEN_1319; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1321 = 12'h529 == io_in ? 12'h3ee : _GEN_1320; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1322 = 12'h52a == io_in ? 12'hb47 : _GEN_1321; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1323 = 12'h52b == io_in ? 12'h3ea : _GEN_1322; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1324 = 12'h52c == io_in ? 12'h408 : _GEN_1323; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1325 = 12'h52d == io_in ? 12'he93 : _GEN_1324; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1326 = 12'h52e == io_in ? 12'hcb : _GEN_1325; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1327 = 12'h52f == io_in ? 12'he31 : _GEN_1326; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1328 = 12'h530 == io_in ? 12'hdcf : _GEN_1327; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1329 = 12'h531 == io_in ? 12'h883 : _GEN_1328; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1330 = 12'h532 == io_in ? 12'h6b1 : _GEN_1329; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1331 = 12'h533 == io_in ? 12'h738 : _GEN_1330; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1332 = 12'h534 == io_in ? 12'h5b2 : _GEN_1331; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1333 = 12'h535 == io_in ? 12'h153 : _GEN_1332; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1334 = 12'h536 == io_in ? 12'hf52 : _GEN_1333; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1335 = 12'h537 == io_in ? 12'hf70 : _GEN_1334; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1336 = 12'h538 == io_in ? 12'hf57 : _GEN_1335; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1337 = 12'h539 == io_in ? 12'hea1 : _GEN_1336; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1338 = 12'h53a == io_in ? 12'he21 : _GEN_1337; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1339 = 12'h53b == io_in ? 12'h1c0 : _GEN_1338; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1340 = 12'h53c == io_in ? 12'h4a0 : _GEN_1339; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1341 = 12'h53d == io_in ? 12'h9ef : _GEN_1340; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1342 = 12'h53e == io_in ? 12'h8ff : _GEN_1341; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1343 = 12'h53f == io_in ? 12'h289 : _GEN_1342; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1344 = 12'h540 == io_in ? 12'he17 : _GEN_1343; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1345 = 12'h541 == io_in ? 12'h4c7 : _GEN_1344; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1346 = 12'h542 == io_in ? 12'hefd : _GEN_1345; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1347 = 12'h543 == io_in ? 12'hb50 : _GEN_1346; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1348 = 12'h544 == io_in ? 12'hc41 : _GEN_1347; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1349 = 12'h545 == io_in ? 12'ha4a : _GEN_1348; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1350 = 12'h546 == io_in ? 12'h85c : _GEN_1349; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1351 = 12'h547 == io_in ? 12'hcbb : _GEN_1350; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1352 = 12'h548 == io_in ? 12'h3db : _GEN_1351; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1353 = 12'h549 == io_in ? 12'ha9d : _GEN_1352; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1354 = 12'h54a == io_in ? 12'hce9 : _GEN_1353; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1355 = 12'h54b == io_in ? 12'hc0f : _GEN_1354; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1356 = 12'h54c == io_in ? 12'h5c6 : _GEN_1355; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1357 = 12'h54d == io_in ? 12'ha49 : _GEN_1356; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1358 = 12'h54e == io_in ? 12'hfc8 : _GEN_1357; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1359 = 12'h54f == io_in ? 12'h425 : _GEN_1358; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1360 = 12'h550 == io_in ? 12'h681 : _GEN_1359; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1361 = 12'h551 == io_in ? 12'hf23 : _GEN_1360; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1362 = 12'h552 == io_in ? 12'h519 : _GEN_1361; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1363 = 12'h553 == io_in ? 12'h2fd : _GEN_1362; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1364 = 12'h554 == io_in ? 12'hf80 : _GEN_1363; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1365 = 12'h555 == io_in ? 12'hc8d : _GEN_1364; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1366 = 12'h556 == io_in ? 12'hda9 : _GEN_1365; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1367 = 12'h557 == io_in ? 12'hd66 : _GEN_1366; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1368 = 12'h558 == io_in ? 12'hf93 : _GEN_1367; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1369 = 12'h559 == io_in ? 12'hbe7 : _GEN_1368; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1370 = 12'h55a == io_in ? 12'hbe : _GEN_1369; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1371 = 12'h55b == io_in ? 12'hd51 : _GEN_1370; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1372 = 12'h55c == io_in ? 12'h82 : _GEN_1371; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1373 = 12'h55d == io_in ? 12'hb8c : _GEN_1372; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1374 = 12'h55e == io_in ? 12'h8e8 : _GEN_1373; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1375 = 12'h55f == io_in ? 12'h233 : _GEN_1374; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1376 = 12'h560 == io_in ? 12'ha92 : _GEN_1375; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1377 = 12'h561 == io_in ? 12'h8d6 : _GEN_1376; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1378 = 12'h562 == io_in ? 12'hf5e : _GEN_1377; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1379 = 12'h563 == io_in ? 12'h5f4 : _GEN_1378; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1380 = 12'h564 == io_in ? 12'hec9 : _GEN_1379; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1381 = 12'h565 == io_in ? 12'h8e2 : _GEN_1380; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1382 = 12'h566 == io_in ? 12'hcbf : _GEN_1381; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1383 = 12'h567 == io_in ? 12'h54e : _GEN_1382; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1384 = 12'h568 == io_in ? 12'hceb : _GEN_1383; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1385 = 12'h569 == io_in ? 12'h2cc : _GEN_1384; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1386 = 12'h56a == io_in ? 12'h5d1 : _GEN_1385; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1387 = 12'h56b == io_in ? 12'hdab : _GEN_1386; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1388 = 12'h56c == io_in ? 12'h842 : _GEN_1387; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1389 = 12'h56d == io_in ? 12'hd71 : _GEN_1388; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1390 = 12'h56e == io_in ? 12'h7cb : _GEN_1389; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1391 = 12'h56f == io_in ? 12'h19b : _GEN_1390; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1392 = 12'h570 == io_in ? 12'hfcd : _GEN_1391; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1393 = 12'h571 == io_in ? 12'he31 : _GEN_1392; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1394 = 12'h572 == io_in ? 12'h8e6 : _GEN_1393; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1395 = 12'h573 == io_in ? 12'ha2b : _GEN_1394; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1396 = 12'h574 == io_in ? 12'h35d : _GEN_1395; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1397 = 12'h575 == io_in ? 12'h66e : _GEN_1396; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1398 = 12'h576 == io_in ? 12'he17 : _GEN_1397; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1399 = 12'h577 == io_in ? 12'h84f : _GEN_1398; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1400 = 12'h578 == io_in ? 12'hbc2 : _GEN_1399; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1401 = 12'h579 == io_in ? 12'he92 : _GEN_1400; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1402 = 12'h57a == io_in ? 12'hb7a : _GEN_1401; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1403 = 12'h57b == io_in ? 12'hcbd : _GEN_1402; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1404 = 12'h57c == io_in ? 12'haeb : _GEN_1403; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1405 = 12'h57d == io_in ? 12'h154 : _GEN_1404; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1406 = 12'h57e == io_in ? 12'h7bd : _GEN_1405; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1407 = 12'h57f == io_in ? 12'h47f : _GEN_1406; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1408 = 12'h580 == io_in ? 12'h2e : _GEN_1407; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1409 = 12'h581 == io_in ? 12'hc54 : _GEN_1408; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1410 = 12'h582 == io_in ? 12'hf44 : _GEN_1409; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1411 = 12'h583 == io_in ? 12'h7a9 : _GEN_1410; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1412 = 12'h584 == io_in ? 12'h264 : _GEN_1411; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1413 = 12'h585 == io_in ? 12'h700 : _GEN_1412; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1414 = 12'h586 == io_in ? 12'he78 : _GEN_1413; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1415 = 12'h587 == io_in ? 12'h988 : _GEN_1414; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1416 = 12'h588 == io_in ? 12'hd74 : _GEN_1415; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1417 = 12'h589 == io_in ? 12'h233 : _GEN_1416; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1418 = 12'h58a == io_in ? 12'h540 : _GEN_1417; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1419 = 12'h58b == io_in ? 12'h517 : _GEN_1418; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1420 = 12'h58c == io_in ? 12'h3aa : _GEN_1419; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1421 = 12'h58d == io_in ? 12'hd48 : _GEN_1420; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1422 = 12'h58e == io_in ? 12'h36c : _GEN_1421; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1423 = 12'h58f == io_in ? 12'hd29 : _GEN_1422; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1424 = 12'h590 == io_in ? 12'h7d5 : _GEN_1423; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1425 = 12'h591 == io_in ? 12'hd75 : _GEN_1424; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1426 = 12'h592 == io_in ? 12'hf19 : _GEN_1425; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1427 = 12'h593 == io_in ? 12'h1b8 : _GEN_1426; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1428 = 12'h594 == io_in ? 12'h5e1 : _GEN_1427; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1429 = 12'h595 == io_in ? 12'h5a6 : _GEN_1428; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1430 = 12'h596 == io_in ? 12'hc1c : _GEN_1429; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1431 = 12'h597 == io_in ? 12'h64c : _GEN_1430; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1432 = 12'h598 == io_in ? 12'hab6 : _GEN_1431; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1433 = 12'h599 == io_in ? 12'hd45 : _GEN_1432; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1434 = 12'h59a == io_in ? 12'hdb4 : _GEN_1433; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1435 = 12'h59b == io_in ? 12'h1d2 : _GEN_1434; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1436 = 12'h59c == io_in ? 12'h5d1 : _GEN_1435; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1437 = 12'h59d == io_in ? 12'h76e : _GEN_1436; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1438 = 12'h59e == io_in ? 12'h98f : _GEN_1437; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1439 = 12'h59f == io_in ? 12'hde1 : _GEN_1438; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1440 = 12'h5a0 == io_in ? 12'h832 : _GEN_1439; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1441 = 12'h5a1 == io_in ? 12'hfe8 : _GEN_1440; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1442 = 12'h5a2 == io_in ? 12'ha5e : _GEN_1441; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1443 = 12'h5a3 == io_in ? 12'h1a : _GEN_1442; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1444 = 12'h5a4 == io_in ? 12'hbcd : _GEN_1443; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1445 = 12'h5a5 == io_in ? 12'h493 : _GEN_1444; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1446 = 12'h5a6 == io_in ? 12'hf41 : _GEN_1445; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1447 = 12'h5a7 == io_in ? 12'h4b : _GEN_1446; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1448 = 12'h5a8 == io_in ? 12'h7a6 : _GEN_1447; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1449 = 12'h5a9 == io_in ? 12'hf16 : _GEN_1448; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1450 = 12'h5aa == io_in ? 12'hfe1 : _GEN_1449; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1451 = 12'h5ab == io_in ? 12'h2fb : _GEN_1450; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1452 = 12'h5ac == io_in ? 12'h909 : _GEN_1451; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1453 = 12'h5ad == io_in ? 12'ha9 : _GEN_1452; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1454 = 12'h5ae == io_in ? 12'h70 : _GEN_1453; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1455 = 12'h5af == io_in ? 12'hb50 : _GEN_1454; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1456 = 12'h5b0 == io_in ? 12'hefb : _GEN_1455; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1457 = 12'h5b1 == io_in ? 12'hfd8 : _GEN_1456; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1458 = 12'h5b2 == io_in ? 12'h730 : _GEN_1457; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1459 = 12'h5b3 == io_in ? 12'h6bf : _GEN_1458; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1460 = 12'h5b4 == io_in ? 12'heb6 : _GEN_1459; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1461 = 12'h5b5 == io_in ? 12'h369 : _GEN_1460; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1462 = 12'h5b6 == io_in ? 12'ha26 : _GEN_1461; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1463 = 12'h5b7 == io_in ? 12'he8e : _GEN_1462; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1464 = 12'h5b8 == io_in ? 12'he43 : _GEN_1463; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1465 = 12'h5b9 == io_in ? 12'he10 : _GEN_1464; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1466 = 12'h5ba == io_in ? 12'h1f : _GEN_1465; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1467 = 12'h5bb == io_in ? 12'h13e : _GEN_1466; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1468 = 12'h5bc == io_in ? 12'h439 : _GEN_1467; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1469 = 12'h5bd == io_in ? 12'h9c0 : _GEN_1468; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1470 = 12'h5be == io_in ? 12'he37 : _GEN_1469; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1471 = 12'h5bf == io_in ? 12'haf3 : _GEN_1470; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1472 = 12'h5c0 == io_in ? 12'h34b : _GEN_1471; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1473 = 12'h5c1 == io_in ? 12'hfd3 : _GEN_1472; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1474 = 12'h5c2 == io_in ? 12'h9e9 : _GEN_1473; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1475 = 12'h5c3 == io_in ? 12'he92 : _GEN_1474; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1476 = 12'h5c4 == io_in ? 12'hf3c : _GEN_1475; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1477 = 12'h5c5 == io_in ? 12'haed : _GEN_1476; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1478 = 12'h5c6 == io_in ? 12'h1f : _GEN_1477; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1479 = 12'h5c7 == io_in ? 12'hc6 : _GEN_1478; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1480 = 12'h5c8 == io_in ? 12'hbb9 : _GEN_1479; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1481 = 12'h5c9 == io_in ? 12'h171 : _GEN_1480; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1482 = 12'h5ca == io_in ? 12'h12f : _GEN_1481; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1483 = 12'h5cb == io_in ? 12'h57b : _GEN_1482; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1484 = 12'h5cc == io_in ? 12'h860 : _GEN_1483; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1485 = 12'h5cd == io_in ? 12'h1f5 : _GEN_1484; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1486 = 12'h5ce == io_in ? 12'hfc6 : _GEN_1485; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1487 = 12'h5cf == io_in ? 12'hb36 : _GEN_1486; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1488 = 12'h5d0 == io_in ? 12'hf25 : _GEN_1487; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1489 = 12'h5d1 == io_in ? 12'h36 : _GEN_1488; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1490 = 12'h5d2 == io_in ? 12'h15f : _GEN_1489; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1491 = 12'h5d3 == io_in ? 12'h5f5 : _GEN_1490; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1492 = 12'h5d4 == io_in ? 12'h9a4 : _GEN_1491; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1493 = 12'h5d5 == io_in ? 12'hf4a : _GEN_1492; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1494 = 12'h5d6 == io_in ? 12'h7a3 : _GEN_1493; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1495 = 12'h5d7 == io_in ? 12'h494 : _GEN_1494; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1496 = 12'h5d8 == io_in ? 12'hbc : _GEN_1495; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1497 = 12'h5d9 == io_in ? 12'hf6c : _GEN_1496; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1498 = 12'h5da == io_in ? 12'h64c : _GEN_1497; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1499 = 12'h5db == io_in ? 12'hcc6 : _GEN_1498; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1500 = 12'h5dc == io_in ? 12'hbe : _GEN_1499; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1501 = 12'h5dd == io_in ? 12'h229 : _GEN_1500; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1502 = 12'h5de == io_in ? 12'hbf1 : _GEN_1501; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1503 = 12'h5df == io_in ? 12'h6bc : _GEN_1502; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1504 = 12'h5e0 == io_in ? 12'hfbf : _GEN_1503; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1505 = 12'h5e1 == io_in ? 12'h985 : _GEN_1504; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1506 = 12'h5e2 == io_in ? 12'h10 : _GEN_1505; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1507 = 12'h5e3 == io_in ? 12'h36f : _GEN_1506; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1508 = 12'h5e4 == io_in ? 12'h6e4 : _GEN_1507; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1509 = 12'h5e5 == io_in ? 12'hdda : _GEN_1508; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1510 = 12'h5e6 == io_in ? 12'hf21 : _GEN_1509; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1511 = 12'h5e7 == io_in ? 12'h3f : _GEN_1510; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1512 = 12'h5e8 == io_in ? 12'h94f : _GEN_1511; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1513 = 12'h5e9 == io_in ? 12'h5ba : _GEN_1512; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1514 = 12'h5ea == io_in ? 12'h729 : _GEN_1513; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1515 = 12'h5eb == io_in ? 12'h56c : _GEN_1514; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1516 = 12'h5ec == io_in ? 12'h197 : _GEN_1515; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1517 = 12'h5ed == io_in ? 12'hb99 : _GEN_1516; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1518 = 12'h5ee == io_in ? 12'h4da : _GEN_1517; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1519 = 12'h5ef == io_in ? 12'h875 : _GEN_1518; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1520 = 12'h5f0 == io_in ? 12'had5 : _GEN_1519; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1521 = 12'h5f1 == io_in ? 12'h1c1 : _GEN_1520; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1522 = 12'h5f2 == io_in ? 12'h115 : _GEN_1521; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1523 = 12'h5f3 == io_in ? 12'h926 : _GEN_1522; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1524 = 12'h5f4 == io_in ? 12'hc74 : _GEN_1523; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1525 = 12'h5f5 == io_in ? 12'hf9a : _GEN_1524; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1526 = 12'h5f6 == io_in ? 12'h63 : _GEN_1525; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1527 = 12'h5f7 == io_in ? 12'ha82 : _GEN_1526; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1528 = 12'h5f8 == io_in ? 12'h43e : _GEN_1527; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1529 = 12'h5f9 == io_in ? 12'h6bd : _GEN_1528; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1530 = 12'h5fa == io_in ? 12'he87 : _GEN_1529; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1531 = 12'h5fb == io_in ? 12'h586 : _GEN_1530; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1532 = 12'h5fc == io_in ? 12'h2e4 : _GEN_1531; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1533 = 12'h5fd == io_in ? 12'h546 : _GEN_1532; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1534 = 12'h5fe == io_in ? 12'hd5b : _GEN_1533; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1535 = 12'h5ff == io_in ? 12'ha00 : _GEN_1534; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1536 = 12'h600 == io_in ? 12'hb64 : _GEN_1535; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1537 = 12'h601 == io_in ? 12'h8ce : _GEN_1536; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1538 = 12'h602 == io_in ? 12'hb9d : _GEN_1537; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1539 = 12'h603 == io_in ? 12'hbad : _GEN_1538; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1540 = 12'h604 == io_in ? 12'h231 : _GEN_1539; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1541 = 12'h605 == io_in ? 12'hd4e : _GEN_1540; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1542 = 12'h606 == io_in ? 12'h262 : _GEN_1541; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1543 = 12'h607 == io_in ? 12'haed : _GEN_1542; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1544 = 12'h608 == io_in ? 12'h6a7 : _GEN_1543; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1545 = 12'h609 == io_in ? 12'h92c : _GEN_1544; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1546 = 12'h60a == io_in ? 12'h54 : _GEN_1545; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1547 = 12'h60b == io_in ? 12'hfa8 : _GEN_1546; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1548 = 12'h60c == io_in ? 12'h839 : _GEN_1547; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1549 = 12'h60d == io_in ? 12'h719 : _GEN_1548; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1550 = 12'h60e == io_in ? 12'hc2d : _GEN_1549; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1551 = 12'h60f == io_in ? 12'h9f8 : _GEN_1550; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1552 = 12'h610 == io_in ? 12'hc0d : _GEN_1551; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1553 = 12'h611 == io_in ? 12'hbf5 : _GEN_1552; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1554 = 12'h612 == io_in ? 12'hbd6 : _GEN_1553; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1555 = 12'h613 == io_in ? 12'h2c1 : _GEN_1554; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1556 = 12'h614 == io_in ? 12'h9a1 : _GEN_1555; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1557 = 12'h615 == io_in ? 12'h661 : _GEN_1556; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1558 = 12'h616 == io_in ? 12'hd45 : _GEN_1557; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1559 = 12'h617 == io_in ? 12'h27b : _GEN_1558; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1560 = 12'h618 == io_in ? 12'hbcd : _GEN_1559; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1561 = 12'h619 == io_in ? 12'hc6d : _GEN_1560; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1562 = 12'h61a == io_in ? 12'h804 : _GEN_1561; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1563 = 12'h61b == io_in ? 12'he48 : _GEN_1562; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1564 = 12'h61c == io_in ? 12'hb3e : _GEN_1563; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1565 = 12'h61d == io_in ? 12'h5cc : _GEN_1564; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1566 = 12'h61e == io_in ? 12'hab6 : _GEN_1565; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1567 = 12'h61f == io_in ? 12'hbad : _GEN_1566; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1568 = 12'h620 == io_in ? 12'h978 : _GEN_1567; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1569 = 12'h621 == io_in ? 12'h495 : _GEN_1568; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1570 = 12'h622 == io_in ? 12'hbf9 : _GEN_1569; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1571 = 12'h623 == io_in ? 12'he78 : _GEN_1570; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1572 = 12'h624 == io_in ? 12'h5ed : _GEN_1571; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1573 = 12'h625 == io_in ? 12'hfa3 : _GEN_1572; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1574 = 12'h626 == io_in ? 12'h86a : _GEN_1573; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1575 = 12'h627 == io_in ? 12'hfde : _GEN_1574; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1576 = 12'h628 == io_in ? 12'h5a0 : _GEN_1575; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1577 = 12'h629 == io_in ? 12'h7a4 : _GEN_1576; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1578 = 12'h62a == io_in ? 12'h411 : _GEN_1577; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1579 = 12'h62b == io_in ? 12'h261 : _GEN_1578; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1580 = 12'h62c == io_in ? 12'h1fe : _GEN_1579; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1581 = 12'h62d == io_in ? 12'h6b5 : _GEN_1580; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1582 = 12'h62e == io_in ? 12'h142 : _GEN_1581; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1583 = 12'h62f == io_in ? 12'h5e9 : _GEN_1582; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1584 = 12'h630 == io_in ? 12'hb0b : _GEN_1583; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1585 = 12'h631 == io_in ? 12'ha14 : _GEN_1584; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1586 = 12'h632 == io_in ? 12'hc63 : _GEN_1585; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1587 = 12'h633 == io_in ? 12'hf7c : _GEN_1586; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1588 = 12'h634 == io_in ? 12'h7da : _GEN_1587; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1589 = 12'h635 == io_in ? 12'h2dd : _GEN_1588; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1590 = 12'h636 == io_in ? 12'he42 : _GEN_1589; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1591 = 12'h637 == io_in ? 12'h718 : _GEN_1590; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1592 = 12'h638 == io_in ? 12'h637 : _GEN_1591; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1593 = 12'h639 == io_in ? 12'hd8b : _GEN_1592; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1594 = 12'h63a == io_in ? 12'h758 : _GEN_1593; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1595 = 12'h63b == io_in ? 12'h5e4 : _GEN_1594; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1596 = 12'h63c == io_in ? 12'he62 : _GEN_1595; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1597 = 12'h63d == io_in ? 12'h672 : _GEN_1596; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1598 = 12'h63e == io_in ? 12'h67b : _GEN_1597; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1599 = 12'h63f == io_in ? 12'ha46 : _GEN_1598; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1600 = 12'h640 == io_in ? 12'h439 : _GEN_1599; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1601 = 12'h641 == io_in ? 12'h31f : _GEN_1600; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1602 = 12'h642 == io_in ? 12'hd78 : _GEN_1601; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1603 = 12'h643 == io_in ? 12'h4da : _GEN_1602; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1604 = 12'h644 == io_in ? 12'h51e : _GEN_1603; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1605 = 12'h645 == io_in ? 12'hc62 : _GEN_1604; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1606 = 12'h646 == io_in ? 12'h5d3 : _GEN_1605; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1607 = 12'h647 == io_in ? 12'h7f4 : _GEN_1606; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1608 = 12'h648 == io_in ? 12'he8c : _GEN_1607; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1609 = 12'h649 == io_in ? 12'h315 : _GEN_1608; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1610 = 12'h64a == io_in ? 12'hd3d : _GEN_1609; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1611 = 12'h64b == io_in ? 12'h691 : _GEN_1610; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1612 = 12'h64c == io_in ? 12'h82a : _GEN_1611; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1613 = 12'h64d == io_in ? 12'h197 : _GEN_1612; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1614 = 12'h64e == io_in ? 12'hbe4 : _GEN_1613; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1615 = 12'h64f == io_in ? 12'h2ab : _GEN_1614; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1616 = 12'h650 == io_in ? 12'h4ca : _GEN_1615; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1617 = 12'h651 == io_in ? 12'h641 : _GEN_1616; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1618 = 12'h652 == io_in ? 12'h22e : _GEN_1617; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1619 = 12'h653 == io_in ? 12'h600 : _GEN_1618; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1620 = 12'h654 == io_in ? 12'h64e : _GEN_1619; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1621 = 12'h655 == io_in ? 12'h79a : _GEN_1620; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1622 = 12'h656 == io_in ? 12'h5b4 : _GEN_1621; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1623 = 12'h657 == io_in ? 12'h2e7 : _GEN_1622; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1624 = 12'h658 == io_in ? 12'h2d8 : _GEN_1623; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1625 = 12'h659 == io_in ? 12'hb08 : _GEN_1624; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1626 = 12'h65a == io_in ? 12'h147 : _GEN_1625; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1627 = 12'h65b == io_in ? 12'h1b4 : _GEN_1626; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1628 = 12'h65c == io_in ? 12'h6ac : _GEN_1627; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1629 = 12'h65d == io_in ? 12'h264 : _GEN_1628; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1630 = 12'h65e == io_in ? 12'h543 : _GEN_1629; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1631 = 12'h65f == io_in ? 12'h673 : _GEN_1630; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1632 = 12'h660 == io_in ? 12'h256 : _GEN_1631; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1633 = 12'h661 == io_in ? 12'hdf1 : _GEN_1632; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1634 = 12'h662 == io_in ? 12'h5ff : _GEN_1633; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1635 = 12'h663 == io_in ? 12'h36b : _GEN_1634; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1636 = 12'h664 == io_in ? 12'hac6 : _GEN_1635; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1637 = 12'h665 == io_in ? 12'hfa2 : _GEN_1636; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1638 = 12'h666 == io_in ? 12'h844 : _GEN_1637; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1639 = 12'h667 == io_in ? 12'hfee : _GEN_1638; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1640 = 12'h668 == io_in ? 12'h8d0 : _GEN_1639; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1641 = 12'h669 == io_in ? 12'hc7f : _GEN_1640; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1642 = 12'h66a == io_in ? 12'hf28 : _GEN_1641; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1643 = 12'h66b == io_in ? 12'hd73 : _GEN_1642; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1644 = 12'h66c == io_in ? 12'h3b7 : _GEN_1643; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1645 = 12'h66d == io_in ? 12'ha92 : _GEN_1644; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1646 = 12'h66e == io_in ? 12'hca8 : _GEN_1645; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1647 = 12'h66f == io_in ? 12'hcea : _GEN_1646; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1648 = 12'h670 == io_in ? 12'h95c : _GEN_1647; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1649 = 12'h671 == io_in ? 12'h819 : _GEN_1648; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1650 = 12'h672 == io_in ? 12'h527 : _GEN_1649; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1651 = 12'h673 == io_in ? 12'hca8 : _GEN_1650; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1652 = 12'h674 == io_in ? 12'h5d2 : _GEN_1651; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1653 = 12'h675 == io_in ? 12'hd13 : _GEN_1652; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1654 = 12'h676 == io_in ? 12'hd00 : _GEN_1653; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1655 = 12'h677 == io_in ? 12'hefa : _GEN_1654; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1656 = 12'h678 == io_in ? 12'h81d : _GEN_1655; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1657 = 12'h679 == io_in ? 12'he7a : _GEN_1656; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1658 = 12'h67a == io_in ? 12'h3dd : _GEN_1657; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1659 = 12'h67b == io_in ? 12'h18 : _GEN_1658; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1660 = 12'h67c == io_in ? 12'h4d6 : _GEN_1659; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1661 = 12'h67d == io_in ? 12'h450 : _GEN_1660; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1662 = 12'h67e == io_in ? 12'h8fc : _GEN_1661; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1663 = 12'h67f == io_in ? 12'h68d : _GEN_1662; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1664 = 12'h680 == io_in ? 12'h82e : _GEN_1663; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1665 = 12'h681 == io_in ? 12'hd31 : _GEN_1664; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1666 = 12'h682 == io_in ? 12'h9ed : _GEN_1665; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1667 = 12'h683 == io_in ? 12'he1e : _GEN_1666; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1668 = 12'h684 == io_in ? 12'hc68 : _GEN_1667; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1669 = 12'h685 == io_in ? 12'hdf1 : _GEN_1668; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1670 = 12'h686 == io_in ? 12'h6ba : _GEN_1669; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1671 = 12'h687 == io_in ? 12'hd7b : _GEN_1670; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1672 = 12'h688 == io_in ? 12'h959 : _GEN_1671; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1673 = 12'h689 == io_in ? 12'h681 : _GEN_1672; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1674 = 12'h68a == io_in ? 12'hcd7 : _GEN_1673; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1675 = 12'h68b == io_in ? 12'ha0f : _GEN_1674; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1676 = 12'h68c == io_in ? 12'hc57 : _GEN_1675; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1677 = 12'h68d == io_in ? 12'h975 : _GEN_1676; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1678 = 12'h68e == io_in ? 12'hd4 : _GEN_1677; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1679 = 12'h68f == io_in ? 12'hab8 : _GEN_1678; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1680 = 12'h690 == io_in ? 12'ha10 : _GEN_1679; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1681 = 12'h691 == io_in ? 12'heed : _GEN_1680; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1682 = 12'h692 == io_in ? 12'h5ce : _GEN_1681; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1683 = 12'h693 == io_in ? 12'hd52 : _GEN_1682; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1684 = 12'h694 == io_in ? 12'hecc : _GEN_1683; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1685 = 12'h695 == io_in ? 12'h8e9 : _GEN_1684; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1686 = 12'h696 == io_in ? 12'ha84 : _GEN_1685; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1687 = 12'h697 == io_in ? 12'h8c : _GEN_1686; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1688 = 12'h698 == io_in ? 12'h3e4 : _GEN_1687; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1689 = 12'h699 == io_in ? 12'hc71 : _GEN_1688; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1690 = 12'h69a == io_in ? 12'h5dd : _GEN_1689; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1691 = 12'h69b == io_in ? 12'hb07 : _GEN_1690; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1692 = 12'h69c == io_in ? 12'h75a : _GEN_1691; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1693 = 12'h69d == io_in ? 12'h3fd : _GEN_1692; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1694 = 12'h69e == io_in ? 12'h76d : _GEN_1693; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1695 = 12'h69f == io_in ? 12'hb48 : _GEN_1694; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1696 = 12'h6a0 == io_in ? 12'hcdc : _GEN_1695; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1697 = 12'h6a1 == io_in ? 12'h2a6 : _GEN_1696; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1698 = 12'h6a2 == io_in ? 12'h15e : _GEN_1697; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1699 = 12'h6a3 == io_in ? 12'he15 : _GEN_1698; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1700 = 12'h6a4 == io_in ? 12'hd61 : _GEN_1699; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1701 = 12'h6a5 == io_in ? 12'hd4 : _GEN_1700; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1702 = 12'h6a6 == io_in ? 12'h722 : _GEN_1701; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1703 = 12'h6a7 == io_in ? 12'h76b : _GEN_1702; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1704 = 12'h6a8 == io_in ? 12'hedf : _GEN_1703; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1705 = 12'h6a9 == io_in ? 12'h979 : _GEN_1704; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1706 = 12'h6aa == io_in ? 12'ha98 : _GEN_1705; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1707 = 12'h6ab == io_in ? 12'hed6 : _GEN_1706; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1708 = 12'h6ac == io_in ? 12'h23a : _GEN_1707; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1709 = 12'h6ad == io_in ? 12'hee7 : _GEN_1708; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1710 = 12'h6ae == io_in ? 12'h588 : _GEN_1709; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1711 = 12'h6af == io_in ? 12'h3ba : _GEN_1710; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1712 = 12'h6b0 == io_in ? 12'hf69 : _GEN_1711; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1713 = 12'h6b1 == io_in ? 12'hf7c : _GEN_1712; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1714 = 12'h6b2 == io_in ? 12'h1a0 : _GEN_1713; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1715 = 12'h6b3 == io_in ? 12'hf3f : _GEN_1714; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1716 = 12'h6b4 == io_in ? 12'hbfb : _GEN_1715; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1717 = 12'h6b5 == io_in ? 12'h1a7 : _GEN_1716; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1718 = 12'h6b6 == io_in ? 12'hd6 : _GEN_1717; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1719 = 12'h6b7 == io_in ? 12'hdb0 : _GEN_1718; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1720 = 12'h6b8 == io_in ? 12'hda3 : _GEN_1719; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1721 = 12'h6b9 == io_in ? 12'hc61 : _GEN_1720; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1722 = 12'h6ba == io_in ? 12'h479 : _GEN_1721; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1723 = 12'h6bb == io_in ? 12'h2b4 : _GEN_1722; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1724 = 12'h6bc == io_in ? 12'ha6 : _GEN_1723; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1725 = 12'h6bd == io_in ? 12'h272 : _GEN_1724; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1726 = 12'h6be == io_in ? 12'h40e : _GEN_1725; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1727 = 12'h6bf == io_in ? 12'hd67 : _GEN_1726; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1728 = 12'h6c0 == io_in ? 12'hb1b : _GEN_1727; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1729 = 12'h6c1 == io_in ? 12'hc42 : _GEN_1728; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1730 = 12'h6c2 == io_in ? 12'h5bc : _GEN_1729; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1731 = 12'h6c3 == io_in ? 12'h187 : _GEN_1730; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1732 = 12'h6c4 == io_in ? 12'hb10 : _GEN_1731; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1733 = 12'h6c5 == io_in ? 12'h3cf : _GEN_1732; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1734 = 12'h6c6 == io_in ? 12'h145 : _GEN_1733; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1735 = 12'h6c7 == io_in ? 12'h8e5 : _GEN_1734; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1736 = 12'h6c8 == io_in ? 12'h3f7 : _GEN_1735; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1737 = 12'h6c9 == io_in ? 12'h12b : _GEN_1736; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1738 = 12'h6ca == io_in ? 12'h1e5 : _GEN_1737; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1739 = 12'h6cb == io_in ? 12'h74b : _GEN_1738; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1740 = 12'h6cc == io_in ? 12'haaf : _GEN_1739; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1741 = 12'h6cd == io_in ? 12'hadc : _GEN_1740; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1742 = 12'h6ce == io_in ? 12'h23c : _GEN_1741; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1743 = 12'h6cf == io_in ? 12'h662 : _GEN_1742; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1744 = 12'h6d0 == io_in ? 12'hee1 : _GEN_1743; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1745 = 12'h6d1 == io_in ? 12'hd4f : _GEN_1744; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1746 = 12'h6d2 == io_in ? 12'h3ca : _GEN_1745; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1747 = 12'h6d3 == io_in ? 12'hefd : _GEN_1746; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1748 = 12'h6d4 == io_in ? 12'h200 : _GEN_1747; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1749 = 12'h6d5 == io_in ? 12'h713 : _GEN_1748; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1750 = 12'h6d6 == io_in ? 12'hf5c : _GEN_1749; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1751 = 12'h6d7 == io_in ? 12'h111 : _GEN_1750; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1752 = 12'h6d8 == io_in ? 12'h266 : _GEN_1751; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1753 = 12'h6d9 == io_in ? 12'he13 : _GEN_1752; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1754 = 12'h6da == io_in ? 12'h761 : _GEN_1753; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1755 = 12'h6db == io_in ? 12'h841 : _GEN_1754; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1756 = 12'h6dc == io_in ? 12'h425 : _GEN_1755; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1757 = 12'h6dd == io_in ? 12'hcac : _GEN_1756; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1758 = 12'h6de == io_in ? 12'h52c : _GEN_1757; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1759 = 12'h6df == io_in ? 12'hc83 : _GEN_1758; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1760 = 12'h6e0 == io_in ? 12'h5ee : _GEN_1759; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1761 = 12'h6e1 == io_in ? 12'h639 : _GEN_1760; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1762 = 12'h6e2 == io_in ? 12'hf9a : _GEN_1761; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1763 = 12'h6e3 == io_in ? 12'hdbc : _GEN_1762; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1764 = 12'h6e4 == io_in ? 12'h9d3 : _GEN_1763; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1765 = 12'h6e5 == io_in ? 12'ha05 : _GEN_1764; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1766 = 12'h6e6 == io_in ? 12'h6fb : _GEN_1765; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1767 = 12'h6e7 == io_in ? 12'h7af : _GEN_1766; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1768 = 12'h6e8 == io_in ? 12'hef5 : _GEN_1767; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1769 = 12'h6e9 == io_in ? 12'hc09 : _GEN_1768; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1770 = 12'h6ea == io_in ? 12'hf9a : _GEN_1769; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1771 = 12'h6eb == io_in ? 12'h5bf : _GEN_1770; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1772 = 12'h6ec == io_in ? 12'h790 : _GEN_1771; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1773 = 12'h6ed == io_in ? 12'hd91 : _GEN_1772; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1774 = 12'h6ee == io_in ? 12'h28f : _GEN_1773; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1775 = 12'h6ef == io_in ? 12'h241 : _GEN_1774; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1776 = 12'h6f0 == io_in ? 12'h885 : _GEN_1775; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1777 = 12'h6f1 == io_in ? 12'h792 : _GEN_1776; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1778 = 12'h6f2 == io_in ? 12'ha33 : _GEN_1777; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1779 = 12'h6f3 == io_in ? 12'hc6b : _GEN_1778; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1780 = 12'h6f4 == io_in ? 12'hbc3 : _GEN_1779; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1781 = 12'h6f5 == io_in ? 12'h716 : _GEN_1780; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1782 = 12'h6f6 == io_in ? 12'hc29 : _GEN_1781; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1783 = 12'h6f7 == io_in ? 12'h4c5 : _GEN_1782; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1784 = 12'h6f8 == io_in ? 12'h295 : _GEN_1783; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1785 = 12'h6f9 == io_in ? 12'h4b1 : _GEN_1784; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1786 = 12'h6fa == io_in ? 12'h31b : _GEN_1785; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1787 = 12'h6fb == io_in ? 12'h83 : _GEN_1786; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1788 = 12'h6fc == io_in ? 12'h20f : _GEN_1787; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1789 = 12'h6fd == io_in ? 12'hced : _GEN_1788; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1790 = 12'h6fe == io_in ? 12'hc5f : _GEN_1789; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1791 = 12'h6ff == io_in ? 12'h6da : _GEN_1790; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1792 = 12'h700 == io_in ? 12'h923 : _GEN_1791; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1793 = 12'h701 == io_in ? 12'h4ae : _GEN_1792; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1794 = 12'h702 == io_in ? 12'hce9 : _GEN_1793; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1795 = 12'h703 == io_in ? 12'hb0e : _GEN_1794; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1796 = 12'h704 == io_in ? 12'haca : _GEN_1795; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1797 = 12'h705 == io_in ? 12'h460 : _GEN_1796; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1798 = 12'h706 == io_in ? 12'h9bd : _GEN_1797; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1799 = 12'h707 == io_in ? 12'h587 : _GEN_1798; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1800 = 12'h708 == io_in ? 12'h79d : _GEN_1799; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1801 = 12'h709 == io_in ? 12'h3f8 : _GEN_1800; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1802 = 12'h70a == io_in ? 12'h475 : _GEN_1801; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1803 = 12'h70b == io_in ? 12'hd1c : _GEN_1802; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1804 = 12'h70c == io_in ? 12'h17b : _GEN_1803; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1805 = 12'h70d == io_in ? 12'hb1e : _GEN_1804; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1806 = 12'h70e == io_in ? 12'h764 : _GEN_1805; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1807 = 12'h70f == io_in ? 12'hf60 : _GEN_1806; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1808 = 12'h710 == io_in ? 12'h459 : _GEN_1807; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1809 = 12'h711 == io_in ? 12'h18c : _GEN_1808; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1810 = 12'h712 == io_in ? 12'h6d3 : _GEN_1809; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1811 = 12'h713 == io_in ? 12'h6c6 : _GEN_1810; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1812 = 12'h714 == io_in ? 12'h3a3 : _GEN_1811; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1813 = 12'h715 == io_in ? 12'h72c : _GEN_1812; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1814 = 12'h716 == io_in ? 12'hf30 : _GEN_1813; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1815 = 12'h717 == io_in ? 12'hc2e : _GEN_1814; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1816 = 12'h718 == io_in ? 12'h994 : _GEN_1815; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1817 = 12'h719 == io_in ? 12'hf54 : _GEN_1816; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1818 = 12'h71a == io_in ? 12'h1b4 : _GEN_1817; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1819 = 12'h71b == io_in ? 12'h6d0 : _GEN_1818; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1820 = 12'h71c == io_in ? 12'ha0e : _GEN_1819; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1821 = 12'h71d == io_in ? 12'h28d : _GEN_1820; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1822 = 12'h71e == io_in ? 12'ha50 : _GEN_1821; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1823 = 12'h71f == io_in ? 12'h23c : _GEN_1822; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1824 = 12'h720 == io_in ? 12'hda2 : _GEN_1823; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1825 = 12'h721 == io_in ? 12'hcea : _GEN_1824; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1826 = 12'h722 == io_in ? 12'h774 : _GEN_1825; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1827 = 12'h723 == io_in ? 12'h305 : _GEN_1826; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1828 = 12'h724 == io_in ? 12'h272 : _GEN_1827; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1829 = 12'h725 == io_in ? 12'h51 : _GEN_1828; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1830 = 12'h726 == io_in ? 12'h57a : _GEN_1829; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1831 = 12'h727 == io_in ? 12'h48e : _GEN_1830; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1832 = 12'h728 == io_in ? 12'haab : _GEN_1831; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1833 = 12'h729 == io_in ? 12'h8b4 : _GEN_1832; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1834 = 12'h72a == io_in ? 12'hfec : _GEN_1833; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1835 = 12'h72b == io_in ? 12'hec2 : _GEN_1834; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1836 = 12'h72c == io_in ? 12'hce6 : _GEN_1835; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1837 = 12'h72d == io_in ? 12'h997 : _GEN_1836; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1838 = 12'h72e == io_in ? 12'h74e : _GEN_1837; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1839 = 12'h72f == io_in ? 12'hab2 : _GEN_1838; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1840 = 12'h730 == io_in ? 12'h78e : _GEN_1839; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1841 = 12'h731 == io_in ? 12'he9d : _GEN_1840; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1842 = 12'h732 == io_in ? 12'h55d : _GEN_1841; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1843 = 12'h733 == io_in ? 12'hecb : _GEN_1842; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1844 = 12'h734 == io_in ? 12'h176 : _GEN_1843; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1845 = 12'h735 == io_in ? 12'ha6d : _GEN_1844; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1846 = 12'h736 == io_in ? 12'h6c5 : _GEN_1845; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1847 = 12'h737 == io_in ? 12'h4ec : _GEN_1846; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1848 = 12'h738 == io_in ? 12'h729 : _GEN_1847; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1849 = 12'h739 == io_in ? 12'h735 : _GEN_1848; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1850 = 12'h73a == io_in ? 12'h9b3 : _GEN_1849; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1851 = 12'h73b == io_in ? 12'h7ea : _GEN_1850; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1852 = 12'h73c == io_in ? 12'hcb7 : _GEN_1851; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1853 = 12'h73d == io_in ? 12'h865 : _GEN_1852; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1854 = 12'h73e == io_in ? 12'h5cd : _GEN_1853; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1855 = 12'h73f == io_in ? 12'hdfc : _GEN_1854; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1856 = 12'h740 == io_in ? 12'h987 : _GEN_1855; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1857 = 12'h741 == io_in ? 12'h62b : _GEN_1856; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1858 = 12'h742 == io_in ? 12'h3b0 : _GEN_1857; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1859 = 12'h743 == io_in ? 12'h87d : _GEN_1858; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1860 = 12'h744 == io_in ? 12'h80d : _GEN_1859; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1861 = 12'h745 == io_in ? 12'h71a : _GEN_1860; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1862 = 12'h746 == io_in ? 12'h8c0 : _GEN_1861; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1863 = 12'h747 == io_in ? 12'h6c1 : _GEN_1862; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1864 = 12'h748 == io_in ? 12'h320 : _GEN_1863; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1865 = 12'h749 == io_in ? 12'h3ba : _GEN_1864; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1866 = 12'h74a == io_in ? 12'hd50 : _GEN_1865; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1867 = 12'h74b == io_in ? 12'h46f : _GEN_1866; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1868 = 12'h74c == io_in ? 12'h1f4 : _GEN_1867; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1869 = 12'h74d == io_in ? 12'h1b9 : _GEN_1868; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1870 = 12'h74e == io_in ? 12'h653 : _GEN_1869; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1871 = 12'h74f == io_in ? 12'hf8a : _GEN_1870; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1872 = 12'h750 == io_in ? 12'h98a : _GEN_1871; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1873 = 12'h751 == io_in ? 12'h9d3 : _GEN_1872; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1874 = 12'h752 == io_in ? 12'hd32 : _GEN_1873; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1875 = 12'h753 == io_in ? 12'h6e1 : _GEN_1874; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1876 = 12'h754 == io_in ? 12'h559 : _GEN_1875; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1877 = 12'h755 == io_in ? 12'hc1c : _GEN_1876; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1878 = 12'h756 == io_in ? 12'hd6e : _GEN_1877; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1879 = 12'h757 == io_in ? 12'h6db : _GEN_1878; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1880 = 12'h758 == io_in ? 12'h2b9 : _GEN_1879; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1881 = 12'h759 == io_in ? 12'hb59 : _GEN_1880; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1882 = 12'h75a == io_in ? 12'hb70 : _GEN_1881; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1883 = 12'h75b == io_in ? 12'hced : _GEN_1882; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1884 = 12'h75c == io_in ? 12'h3c9 : _GEN_1883; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1885 = 12'h75d == io_in ? 12'h1c9 : _GEN_1884; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1886 = 12'h75e == io_in ? 12'he33 : _GEN_1885; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1887 = 12'h75f == io_in ? 12'h5f4 : _GEN_1886; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1888 = 12'h760 == io_in ? 12'h417 : _GEN_1887; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1889 = 12'h761 == io_in ? 12'h9f9 : _GEN_1888; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1890 = 12'h762 == io_in ? 12'hfdd : _GEN_1889; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1891 = 12'h763 == io_in ? 12'h1d9 : _GEN_1890; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1892 = 12'h764 == io_in ? 12'h5dd : _GEN_1891; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1893 = 12'h765 == io_in ? 12'h5aa : _GEN_1892; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1894 = 12'h766 == io_in ? 12'h236 : _GEN_1893; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1895 = 12'h767 == io_in ? 12'h81 : _GEN_1894; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1896 = 12'h768 == io_in ? 12'h168 : _GEN_1895; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1897 = 12'h769 == io_in ? 12'hdcb : _GEN_1896; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1898 = 12'h76a == io_in ? 12'hb41 : _GEN_1897; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1899 = 12'h76b == io_in ? 12'he3d : _GEN_1898; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1900 = 12'h76c == io_in ? 12'hf26 : _GEN_1899; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1901 = 12'h76d == io_in ? 12'ha2f : _GEN_1900; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1902 = 12'h76e == io_in ? 12'hcf1 : _GEN_1901; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1903 = 12'h76f == io_in ? 12'h630 : _GEN_1902; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1904 = 12'h770 == io_in ? 12'hbd : _GEN_1903; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1905 = 12'h771 == io_in ? 12'h10e : _GEN_1904; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1906 = 12'h772 == io_in ? 12'h7ab : _GEN_1905; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1907 = 12'h773 == io_in ? 12'h95c : _GEN_1906; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1908 = 12'h774 == io_in ? 12'h754 : _GEN_1907; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1909 = 12'h775 == io_in ? 12'h6d1 : _GEN_1908; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1910 = 12'h776 == io_in ? 12'h909 : _GEN_1909; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1911 = 12'h777 == io_in ? 12'hb25 : _GEN_1910; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1912 = 12'h778 == io_in ? 12'h53 : _GEN_1911; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1913 = 12'h779 == io_in ? 12'h1dd : _GEN_1912; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1914 = 12'h77a == io_in ? 12'hca5 : _GEN_1913; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1915 = 12'h77b == io_in ? 12'he51 : _GEN_1914; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1916 = 12'h77c == io_in ? 12'h944 : _GEN_1915; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1917 = 12'h77d == io_in ? 12'h60c : _GEN_1916; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1918 = 12'h77e == io_in ? 12'h11e : _GEN_1917; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1919 = 12'h77f == io_in ? 12'he9e : _GEN_1918; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1920 = 12'h780 == io_in ? 12'h579 : _GEN_1919; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1921 = 12'h781 == io_in ? 12'hc12 : _GEN_1920; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1922 = 12'h782 == io_in ? 12'hb75 : _GEN_1921; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1923 = 12'h783 == io_in ? 12'hd51 : _GEN_1922; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1924 = 12'h784 == io_in ? 12'h229 : _GEN_1923; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1925 = 12'h785 == io_in ? 12'h50c : _GEN_1924; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1926 = 12'h786 == io_in ? 12'hb6a : _GEN_1925; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1927 = 12'h787 == io_in ? 12'h62c : _GEN_1926; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1928 = 12'h788 == io_in ? 12'h84a : _GEN_1927; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1929 = 12'h789 == io_in ? 12'hdf7 : _GEN_1928; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1930 = 12'h78a == io_in ? 12'h571 : _GEN_1929; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1931 = 12'h78b == io_in ? 12'hcaa : _GEN_1930; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1932 = 12'h78c == io_in ? 12'hed6 : _GEN_1931; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1933 = 12'h78d == io_in ? 12'h55c : _GEN_1932; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1934 = 12'h78e == io_in ? 12'h684 : _GEN_1933; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1935 = 12'h78f == io_in ? 12'hf77 : _GEN_1934; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1936 = 12'h790 == io_in ? 12'hf4a : _GEN_1935; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1937 = 12'h791 == io_in ? 12'hbab : _GEN_1936; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1938 = 12'h792 == io_in ? 12'h2b3 : _GEN_1937; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1939 = 12'h793 == io_in ? 12'hccc : _GEN_1938; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1940 = 12'h794 == io_in ? 12'h3c5 : _GEN_1939; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1941 = 12'h795 == io_in ? 12'h26 : _GEN_1940; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1942 = 12'h796 == io_in ? 12'hb36 : _GEN_1941; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1943 = 12'h797 == io_in ? 12'h267 : _GEN_1942; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1944 = 12'h798 == io_in ? 12'hf8a : _GEN_1943; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1945 = 12'h799 == io_in ? 12'h6ca : _GEN_1944; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1946 = 12'h79a == io_in ? 12'ha61 : _GEN_1945; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1947 = 12'h79b == io_in ? 12'h703 : _GEN_1946; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1948 = 12'h79c == io_in ? 12'h550 : _GEN_1947; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1949 = 12'h79d == io_in ? 12'h29b : _GEN_1948; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1950 = 12'h79e == io_in ? 12'hb71 : _GEN_1949; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1951 = 12'h79f == io_in ? 12'h234 : _GEN_1950; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1952 = 12'h7a0 == io_in ? 12'ha48 : _GEN_1951; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1953 = 12'h7a1 == io_in ? 12'h1e8 : _GEN_1952; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1954 = 12'h7a2 == io_in ? 12'heed : _GEN_1953; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1955 = 12'h7a3 == io_in ? 12'h745 : _GEN_1954; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1956 = 12'h7a4 == io_in ? 12'h919 : _GEN_1955; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1957 = 12'h7a5 == io_in ? 12'hb5f : _GEN_1956; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1958 = 12'h7a6 == io_in ? 12'h8e4 : _GEN_1957; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1959 = 12'h7a7 == io_in ? 12'hcc7 : _GEN_1958; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1960 = 12'h7a8 == io_in ? 12'h7af : _GEN_1959; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1961 = 12'h7a9 == io_in ? 12'ha38 : _GEN_1960; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1962 = 12'h7aa == io_in ? 12'h8b8 : _GEN_1961; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1963 = 12'h7ab == io_in ? 12'heb7 : _GEN_1962; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1964 = 12'h7ac == io_in ? 12'h784 : _GEN_1963; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1965 = 12'h7ad == io_in ? 12'h9c1 : _GEN_1964; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1966 = 12'h7ae == io_in ? 12'heee : _GEN_1965; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1967 = 12'h7af == io_in ? 12'h570 : _GEN_1966; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1968 = 12'h7b0 == io_in ? 12'h77d : _GEN_1967; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1969 = 12'h7b1 == io_in ? 12'h4cd : _GEN_1968; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1970 = 12'h7b2 == io_in ? 12'h7ab : _GEN_1969; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1971 = 12'h7b3 == io_in ? 12'he59 : _GEN_1970; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1972 = 12'h7b4 == io_in ? 12'hca6 : _GEN_1971; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1973 = 12'h7b5 == io_in ? 12'h102 : _GEN_1972; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1974 = 12'h7b6 == io_in ? 12'hb21 : _GEN_1973; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1975 = 12'h7b7 == io_in ? 12'h1de : _GEN_1974; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1976 = 12'h7b8 == io_in ? 12'hc1d : _GEN_1975; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1977 = 12'h7b9 == io_in ? 12'h7b : _GEN_1976; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1978 = 12'h7ba == io_in ? 12'h93e : _GEN_1977; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1979 = 12'h7bb == io_in ? 12'hf81 : _GEN_1978; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1980 = 12'h7bc == io_in ? 12'haed : _GEN_1979; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1981 = 12'h7bd == io_in ? 12'hba7 : _GEN_1980; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1982 = 12'h7be == io_in ? 12'hdae : _GEN_1981; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1983 = 12'h7bf == io_in ? 12'h6eb : _GEN_1982; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1984 = 12'h7c0 == io_in ? 12'h2f0 : _GEN_1983; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1985 = 12'h7c1 == io_in ? 12'h1a3 : _GEN_1984; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1986 = 12'h7c2 == io_in ? 12'hbbf : _GEN_1985; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1987 = 12'h7c3 == io_in ? 12'haa2 : _GEN_1986; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1988 = 12'h7c4 == io_in ? 12'hf5c : _GEN_1987; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1989 = 12'h7c5 == io_in ? 12'hd63 : _GEN_1988; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1990 = 12'h7c6 == io_in ? 12'h794 : _GEN_1989; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1991 = 12'h7c7 == io_in ? 12'h5b8 : _GEN_1990; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1992 = 12'h7c8 == io_in ? 12'hd2e : _GEN_1991; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1993 = 12'h7c9 == io_in ? 12'h1a9 : _GEN_1992; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1994 = 12'h7ca == io_in ? 12'h978 : _GEN_1993; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1995 = 12'h7cb == io_in ? 12'hc10 : _GEN_1994; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1996 = 12'h7cc == io_in ? 12'hef4 : _GEN_1995; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1997 = 12'h7cd == io_in ? 12'hce9 : _GEN_1996; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1998 = 12'h7ce == io_in ? 12'h797 : _GEN_1997; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_1999 = 12'h7cf == io_in ? 12'h923 : _GEN_1998; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2000 = 12'h7d0 == io_in ? 12'he : _GEN_1999; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2001 = 12'h7d1 == io_in ? 12'h12c : _GEN_2000; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2002 = 12'h7d2 == io_in ? 12'hea3 : _GEN_2001; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2003 = 12'h7d3 == io_in ? 12'ha37 : _GEN_2002; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2004 = 12'h7d4 == io_in ? 12'h79a : _GEN_2003; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2005 = 12'h7d5 == io_in ? 12'h268 : _GEN_2004; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2006 = 12'h7d6 == io_in ? 12'h8d : _GEN_2005; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2007 = 12'h7d7 == io_in ? 12'hfa8 : _GEN_2006; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2008 = 12'h7d8 == io_in ? 12'h877 : _GEN_2007; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2009 = 12'h7d9 == io_in ? 12'h196 : _GEN_2008; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2010 = 12'h7da == io_in ? 12'hbf1 : _GEN_2009; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2011 = 12'h7db == io_in ? 12'h913 : _GEN_2010; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2012 = 12'h7dc == io_in ? 12'hb7d : _GEN_2011; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2013 = 12'h7dd == io_in ? 12'h356 : _GEN_2012; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2014 = 12'h7de == io_in ? 12'hb98 : _GEN_2013; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2015 = 12'h7df == io_in ? 12'h632 : _GEN_2014; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2016 = 12'h7e0 == io_in ? 12'h6de : _GEN_2015; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2017 = 12'h7e1 == io_in ? 12'hc3 : _GEN_2016; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2018 = 12'h7e2 == io_in ? 12'hcd2 : _GEN_2017; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2019 = 12'h7e3 == io_in ? 12'h360 : _GEN_2018; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2020 = 12'h7e4 == io_in ? 12'h5a2 : _GEN_2019; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2021 = 12'h7e5 == io_in ? 12'h899 : _GEN_2020; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2022 = 12'h7e6 == io_in ? 12'hf89 : _GEN_2021; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2023 = 12'h7e7 == io_in ? 12'hd8b : _GEN_2022; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2024 = 12'h7e8 == io_in ? 12'h276 : _GEN_2023; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2025 = 12'h7e9 == io_in ? 12'h83a : _GEN_2024; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2026 = 12'h7ea == io_in ? 12'h451 : _GEN_2025; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2027 = 12'h7eb == io_in ? 12'h347 : _GEN_2026; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2028 = 12'h7ec == io_in ? 12'h817 : _GEN_2027; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2029 = 12'h7ed == io_in ? 12'h8ec : _GEN_2028; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2030 = 12'h7ee == io_in ? 12'hbbb : _GEN_2029; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2031 = 12'h7ef == io_in ? 12'h55f : _GEN_2030; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2032 = 12'h7f0 == io_in ? 12'h3d : _GEN_2031; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2033 = 12'h7f1 == io_in ? 12'h879 : _GEN_2032; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2034 = 12'h7f2 == io_in ? 12'h5e1 : _GEN_2033; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2035 = 12'h7f3 == io_in ? 12'ha1f : _GEN_2034; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2036 = 12'h7f4 == io_in ? 12'hd0 : _GEN_2035; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2037 = 12'h7f5 == io_in ? 12'h6de : _GEN_2036; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2038 = 12'h7f6 == io_in ? 12'h83a : _GEN_2037; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2039 = 12'h7f7 == io_in ? 12'h618 : _GEN_2038; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2040 = 12'h7f8 == io_in ? 12'h9f6 : _GEN_2039; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2041 = 12'h7f9 == io_in ? 12'h8d : _GEN_2040; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2042 = 12'h7fa == io_in ? 12'h825 : _GEN_2041; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2043 = 12'h7fb == io_in ? 12'h10c : _GEN_2042; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2044 = 12'h7fc == io_in ? 12'h912 : _GEN_2043; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2045 = 12'h7fd == io_in ? 12'hf93 : _GEN_2044; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2046 = 12'h7fe == io_in ? 12'hf2b : _GEN_2045; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2047 = 12'h7ff == io_in ? 12'hd0e : _GEN_2046; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2048 = 12'h800 == io_in ? 12'h37d : _GEN_2047; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2049 = 12'h801 == io_in ? 12'ha45 : _GEN_2048; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2050 = 12'h802 == io_in ? 12'hf23 : _GEN_2049; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2051 = 12'h803 == io_in ? 12'hb02 : _GEN_2050; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2052 = 12'h804 == io_in ? 12'h4e4 : _GEN_2051; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2053 = 12'h805 == io_in ? 12'hde9 : _GEN_2052; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2054 = 12'h806 == io_in ? 12'h3ff : _GEN_2053; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2055 = 12'h807 == io_in ? 12'h5d0 : _GEN_2054; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2056 = 12'h808 == io_in ? 12'h17b : _GEN_2055; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2057 = 12'h809 == io_in ? 12'hc06 : _GEN_2056; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2058 = 12'h80a == io_in ? 12'h121 : _GEN_2057; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2059 = 12'h80b == io_in ? 12'h423 : _GEN_2058; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2060 = 12'h80c == io_in ? 12'h3cd : _GEN_2059; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2061 = 12'h80d == io_in ? 12'h47d : _GEN_2060; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2062 = 12'h80e == io_in ? 12'hc07 : _GEN_2061; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2063 = 12'h80f == io_in ? 12'he94 : _GEN_2062; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2064 = 12'h810 == io_in ? 12'hbb5 : _GEN_2063; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2065 = 12'h811 == io_in ? 12'ha4d : _GEN_2064; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2066 = 12'h812 == io_in ? 12'h5ba : _GEN_2065; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2067 = 12'h813 == io_in ? 12'h1e6 : _GEN_2066; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2068 = 12'h814 == io_in ? 12'hab2 : _GEN_2067; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2069 = 12'h815 == io_in ? 12'h861 : _GEN_2068; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2070 = 12'h816 == io_in ? 12'h992 : _GEN_2069; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2071 = 12'h817 == io_in ? 12'h615 : _GEN_2070; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2072 = 12'h818 == io_in ? 12'hf04 : _GEN_2071; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2073 = 12'h819 == io_in ? 12'hcb8 : _GEN_2072; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2074 = 12'h81a == io_in ? 12'h1a4 : _GEN_2073; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2075 = 12'h81b == io_in ? 12'h419 : _GEN_2074; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2076 = 12'h81c == io_in ? 12'hf98 : _GEN_2075; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2077 = 12'h81d == io_in ? 12'h661 : _GEN_2076; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2078 = 12'h81e == io_in ? 12'h6de : _GEN_2077; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2079 = 12'h81f == io_in ? 12'hd79 : _GEN_2078; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2080 = 12'h820 == io_in ? 12'hf07 : _GEN_2079; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2081 = 12'h821 == io_in ? 12'h460 : _GEN_2080; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2082 = 12'h822 == io_in ? 12'hac9 : _GEN_2081; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2083 = 12'h823 == io_in ? 12'h732 : _GEN_2082; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2084 = 12'h824 == io_in ? 12'hb7e : _GEN_2083; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2085 = 12'h825 == io_in ? 12'h4e4 : _GEN_2084; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2086 = 12'h826 == io_in ? 12'h8b3 : _GEN_2085; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2087 = 12'h827 == io_in ? 12'h203 : _GEN_2086; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2088 = 12'h828 == io_in ? 12'h67a : _GEN_2087; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2089 = 12'h829 == io_in ? 12'hc2c : _GEN_2088; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2090 = 12'h82a == io_in ? 12'h5d : _GEN_2089; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2091 = 12'h82b == io_in ? 12'hdf5 : _GEN_2090; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2092 = 12'h82c == io_in ? 12'hc6c : _GEN_2091; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2093 = 12'h82d == io_in ? 12'h58a : _GEN_2092; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2094 = 12'h82e == io_in ? 12'h986 : _GEN_2093; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2095 = 12'h82f == io_in ? 12'h7c4 : _GEN_2094; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2096 = 12'h830 == io_in ? 12'h644 : _GEN_2095; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2097 = 12'h831 == io_in ? 12'h6af : _GEN_2096; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2098 = 12'h832 == io_in ? 12'h8b9 : _GEN_2097; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2099 = 12'h833 == io_in ? 12'h215 : _GEN_2098; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2100 = 12'h834 == io_in ? 12'h266 : _GEN_2099; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2101 = 12'h835 == io_in ? 12'h2e8 : _GEN_2100; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2102 = 12'h836 == io_in ? 12'h5b0 : _GEN_2101; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2103 = 12'h837 == io_in ? 12'h8d : _GEN_2102; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2104 = 12'h838 == io_in ? 12'h708 : _GEN_2103; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2105 = 12'h839 == io_in ? 12'h8fb : _GEN_2104; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2106 = 12'h83a == io_in ? 12'h3d4 : _GEN_2105; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2107 = 12'h83b == io_in ? 12'h9ae : _GEN_2106; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2108 = 12'h83c == io_in ? 12'hcca : _GEN_2107; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2109 = 12'h83d == io_in ? 12'h8c8 : _GEN_2108; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2110 = 12'h83e == io_in ? 12'h740 : _GEN_2109; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2111 = 12'h83f == io_in ? 12'h8d9 : _GEN_2110; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2112 = 12'h840 == io_in ? 12'h721 : _GEN_2111; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2113 = 12'h841 == io_in ? 12'hdcf : _GEN_2112; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2114 = 12'h842 == io_in ? 12'h441 : _GEN_2113; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2115 = 12'h843 == io_in ? 12'h264 : _GEN_2114; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2116 = 12'h844 == io_in ? 12'h315 : _GEN_2115; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2117 = 12'h845 == io_in ? 12'hf8d : _GEN_2116; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2118 = 12'h846 == io_in ? 12'h490 : _GEN_2117; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2119 = 12'h847 == io_in ? 12'hf82 : _GEN_2118; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2120 = 12'h848 == io_in ? 12'h7ce : _GEN_2119; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2121 = 12'h849 == io_in ? 12'h941 : _GEN_2120; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2122 = 12'h84a == io_in ? 12'hab1 : _GEN_2121; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2123 = 12'h84b == io_in ? 12'ha0b : _GEN_2122; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2124 = 12'h84c == io_in ? 12'h420 : _GEN_2123; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2125 = 12'h84d == io_in ? 12'h66e : _GEN_2124; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2126 = 12'h84e == io_in ? 12'h7df : _GEN_2125; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2127 = 12'h84f == io_in ? 12'h47c : _GEN_2126; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2128 = 12'h850 == io_in ? 12'h763 : _GEN_2127; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2129 = 12'h851 == io_in ? 12'h222 : _GEN_2128; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2130 = 12'h852 == io_in ? 12'h17 : _GEN_2129; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2131 = 12'h853 == io_in ? 12'h89a : _GEN_2130; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2132 = 12'h854 == io_in ? 12'h120 : _GEN_2131; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2133 = 12'h855 == io_in ? 12'h377 : _GEN_2132; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2134 = 12'h856 == io_in ? 12'h7af : _GEN_2133; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2135 = 12'h857 == io_in ? 12'hef2 : _GEN_2134; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2136 = 12'h858 == io_in ? 12'h419 : _GEN_2135; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2137 = 12'h859 == io_in ? 12'h3f9 : _GEN_2136; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2138 = 12'h85a == io_in ? 12'h185 : _GEN_2137; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2139 = 12'h85b == io_in ? 12'hf6e : _GEN_2138; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2140 = 12'h85c == io_in ? 12'hef0 : _GEN_2139; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2141 = 12'h85d == io_in ? 12'h446 : _GEN_2140; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2142 = 12'h85e == io_in ? 12'h7d5 : _GEN_2141; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2143 = 12'h85f == io_in ? 12'hb87 : _GEN_2142; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2144 = 12'h860 == io_in ? 12'h34a : _GEN_2143; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2145 = 12'h861 == io_in ? 12'haa7 : _GEN_2144; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2146 = 12'h862 == io_in ? 12'he10 : _GEN_2145; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2147 = 12'h863 == io_in ? 12'h692 : _GEN_2146; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2148 = 12'h864 == io_in ? 12'h753 : _GEN_2147; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2149 = 12'h865 == io_in ? 12'h6b4 : _GEN_2148; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2150 = 12'h866 == io_in ? 12'h9a8 : _GEN_2149; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2151 = 12'h867 == io_in ? 12'h9a : _GEN_2150; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2152 = 12'h868 == io_in ? 12'hb90 : _GEN_2151; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2153 = 12'h869 == io_in ? 12'h74b : _GEN_2152; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2154 = 12'h86a == io_in ? 12'haf5 : _GEN_2153; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2155 = 12'h86b == io_in ? 12'ha22 : _GEN_2154; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2156 = 12'h86c == io_in ? 12'he17 : _GEN_2155; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2157 = 12'h86d == io_in ? 12'h5b0 : _GEN_2156; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2158 = 12'h86e == io_in ? 12'hee3 : _GEN_2157; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2159 = 12'h86f == io_in ? 12'hfe5 : _GEN_2158; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2160 = 12'h870 == io_in ? 12'h588 : _GEN_2159; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2161 = 12'h871 == io_in ? 12'hd4b : _GEN_2160; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2162 = 12'h872 == io_in ? 12'hc80 : _GEN_2161; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2163 = 12'h873 == io_in ? 12'h78a : _GEN_2162; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2164 = 12'h874 == io_in ? 12'h241 : _GEN_2163; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2165 = 12'h875 == io_in ? 12'h3c8 : _GEN_2164; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2166 = 12'h876 == io_in ? 12'he4a : _GEN_2165; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2167 = 12'h877 == io_in ? 12'h2d2 : _GEN_2166; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2168 = 12'h878 == io_in ? 12'he8e : _GEN_2167; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2169 = 12'h879 == io_in ? 12'h5e0 : _GEN_2168; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2170 = 12'h87a == io_in ? 12'h308 : _GEN_2169; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2171 = 12'h87b == io_in ? 12'hcb6 : _GEN_2170; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2172 = 12'h87c == io_in ? 12'h27c : _GEN_2171; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2173 = 12'h87d == io_in ? 12'h2de : _GEN_2172; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2174 = 12'h87e == io_in ? 12'h351 : _GEN_2173; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2175 = 12'h87f == io_in ? 12'h162 : _GEN_2174; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2176 = 12'h880 == io_in ? 12'h31b : _GEN_2175; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2177 = 12'h881 == io_in ? 12'h8c7 : _GEN_2176; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2178 = 12'h882 == io_in ? 12'h2b1 : _GEN_2177; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2179 = 12'h883 == io_in ? 12'h1ff : _GEN_2178; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2180 = 12'h884 == io_in ? 12'h56c : _GEN_2179; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2181 = 12'h885 == io_in ? 12'h6e6 : _GEN_2180; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2182 = 12'h886 == io_in ? 12'ha7d : _GEN_2181; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2183 = 12'h887 == io_in ? 12'h29f : _GEN_2182; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2184 = 12'h888 == io_in ? 12'h30b : _GEN_2183; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2185 = 12'h889 == io_in ? 12'h950 : _GEN_2184; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2186 = 12'h88a == io_in ? 12'ha71 : _GEN_2185; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2187 = 12'h88b == io_in ? 12'h2f9 : _GEN_2186; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2188 = 12'h88c == io_in ? 12'ha7e : _GEN_2187; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2189 = 12'h88d == io_in ? 12'h854 : _GEN_2188; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2190 = 12'h88e == io_in ? 12'h36a : _GEN_2189; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2191 = 12'h88f == io_in ? 12'hdf : _GEN_2190; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2192 = 12'h890 == io_in ? 12'h153 : _GEN_2191; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2193 = 12'h891 == io_in ? 12'h821 : _GEN_2192; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2194 = 12'h892 == io_in ? 12'h330 : _GEN_2193; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2195 = 12'h893 == io_in ? 12'h9ed : _GEN_2194; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2196 = 12'h894 == io_in ? 12'h647 : _GEN_2195; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2197 = 12'h895 == io_in ? 12'ha77 : _GEN_2196; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2198 = 12'h896 == io_in ? 12'h6d1 : _GEN_2197; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2199 = 12'h897 == io_in ? 12'h46f : _GEN_2198; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2200 = 12'h898 == io_in ? 12'h257 : _GEN_2199; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2201 = 12'h899 == io_in ? 12'hbb7 : _GEN_2200; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2202 = 12'h89a == io_in ? 12'haa0 : _GEN_2201; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2203 = 12'h89b == io_in ? 12'h62b : _GEN_2202; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2204 = 12'h89c == io_in ? 12'h669 : _GEN_2203; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2205 = 12'h89d == io_in ? 12'h1ad : _GEN_2204; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2206 = 12'h89e == io_in ? 12'h31d : _GEN_2205; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2207 = 12'h89f == io_in ? 12'hb76 : _GEN_2206; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2208 = 12'h8a0 == io_in ? 12'h57 : _GEN_2207; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2209 = 12'h8a1 == io_in ? 12'h3d0 : _GEN_2208; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2210 = 12'h8a2 == io_in ? 12'hed7 : _GEN_2209; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2211 = 12'h8a3 == io_in ? 12'he0f : _GEN_2210; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2212 = 12'h8a4 == io_in ? 12'hc79 : _GEN_2211; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2213 = 12'h8a5 == io_in ? 12'h5e5 : _GEN_2212; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2214 = 12'h8a6 == io_in ? 12'h49d : _GEN_2213; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2215 = 12'h8a7 == io_in ? 12'h712 : _GEN_2214; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2216 = 12'h8a8 == io_in ? 12'h3fe : _GEN_2215; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2217 = 12'h8a9 == io_in ? 12'he77 : _GEN_2216; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2218 = 12'h8aa == io_in ? 12'h76f : _GEN_2217; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2219 = 12'h8ab == io_in ? 12'hae8 : _GEN_2218; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2220 = 12'h8ac == io_in ? 12'hd4c : _GEN_2219; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2221 = 12'h8ad == io_in ? 12'h6ba : _GEN_2220; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2222 = 12'h8ae == io_in ? 12'hf83 : _GEN_2221; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2223 = 12'h8af == io_in ? 12'h32d : _GEN_2222; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2224 = 12'h8b0 == io_in ? 12'h87e : _GEN_2223; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2225 = 12'h8b1 == io_in ? 12'h8ae : _GEN_2224; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2226 = 12'h8b2 == io_in ? 12'h754 : _GEN_2225; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2227 = 12'h8b3 == io_in ? 12'he9f : _GEN_2226; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2228 = 12'h8b4 == io_in ? 12'ha91 : _GEN_2227; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2229 = 12'h8b5 == io_in ? 12'h7d0 : _GEN_2228; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2230 = 12'h8b6 == io_in ? 12'h168 : _GEN_2229; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2231 = 12'h8b7 == io_in ? 12'h87a : _GEN_2230; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2232 = 12'h8b8 == io_in ? 12'he26 : _GEN_2231; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2233 = 12'h8b9 == io_in ? 12'h84c : _GEN_2232; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2234 = 12'h8ba == io_in ? 12'h738 : _GEN_2233; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2235 = 12'h8bb == io_in ? 12'h963 : _GEN_2234; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2236 = 12'h8bc == io_in ? 12'hf73 : _GEN_2235; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2237 = 12'h8bd == io_in ? 12'h611 : _GEN_2236; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2238 = 12'h8be == io_in ? 12'he2a : _GEN_2237; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2239 = 12'h8bf == io_in ? 12'heae : _GEN_2238; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2240 = 12'h8c0 == io_in ? 12'hcc3 : _GEN_2239; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2241 = 12'h8c1 == io_in ? 12'hac : _GEN_2240; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2242 = 12'h8c2 == io_in ? 12'h3fb : _GEN_2241; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2243 = 12'h8c3 == io_in ? 12'h32 : _GEN_2242; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2244 = 12'h8c4 == io_in ? 12'h6a1 : _GEN_2243; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2245 = 12'h8c5 == io_in ? 12'h8b7 : _GEN_2244; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2246 = 12'h8c6 == io_in ? 12'h886 : _GEN_2245; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2247 = 12'h8c7 == io_in ? 12'h7e0 : _GEN_2246; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2248 = 12'h8c8 == io_in ? 12'h7ae : _GEN_2247; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2249 = 12'h8c9 == io_in ? 12'h8af : _GEN_2248; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2250 = 12'h8ca == io_in ? 12'he20 : _GEN_2249; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2251 = 12'h8cb == io_in ? 12'h48b : _GEN_2250; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2252 = 12'h8cc == io_in ? 12'h7e1 : _GEN_2251; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2253 = 12'h8cd == io_in ? 12'hc0d : _GEN_2252; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2254 = 12'h8ce == io_in ? 12'h1ec : _GEN_2253; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2255 = 12'h8cf == io_in ? 12'hdb4 : _GEN_2254; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2256 = 12'h8d0 == io_in ? 12'h8a9 : _GEN_2255; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2257 = 12'h8d1 == io_in ? 12'hd67 : _GEN_2256; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2258 = 12'h8d2 == io_in ? 12'hfc6 : _GEN_2257; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2259 = 12'h8d3 == io_in ? 12'h13d : _GEN_2258; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2260 = 12'h8d4 == io_in ? 12'hdeb : _GEN_2259; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2261 = 12'h8d5 == io_in ? 12'h71b : _GEN_2260; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2262 = 12'h8d6 == io_in ? 12'h69a : _GEN_2261; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2263 = 12'h8d7 == io_in ? 12'h4cd : _GEN_2262; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2264 = 12'h8d8 == io_in ? 12'hc6c : _GEN_2263; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2265 = 12'h8d9 == io_in ? 12'h2a4 : _GEN_2264; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2266 = 12'h8da == io_in ? 12'hd72 : _GEN_2265; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2267 = 12'h8db == io_in ? 12'h892 : _GEN_2266; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2268 = 12'h8dc == io_in ? 12'h217 : _GEN_2267; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2269 = 12'h8dd == io_in ? 12'h964 : _GEN_2268; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2270 = 12'h8de == io_in ? 12'h31b : _GEN_2269; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2271 = 12'h8df == io_in ? 12'h39d : _GEN_2270; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2272 = 12'h8e0 == io_in ? 12'h3de : _GEN_2271; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2273 = 12'h8e1 == io_in ? 12'h8ad : _GEN_2272; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2274 = 12'h8e2 == io_in ? 12'hb3b : _GEN_2273; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2275 = 12'h8e3 == io_in ? 12'hcd3 : _GEN_2274; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2276 = 12'h8e4 == io_in ? 12'h30f : _GEN_2275; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2277 = 12'h8e5 == io_in ? 12'h240 : _GEN_2276; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2278 = 12'h8e6 == io_in ? 12'h6e8 : _GEN_2277; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2279 = 12'h8e7 == io_in ? 12'hea6 : _GEN_2278; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2280 = 12'h8e8 == io_in ? 12'h7ca : _GEN_2279; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2281 = 12'h8e9 == io_in ? 12'h4f7 : _GEN_2280; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2282 = 12'h8ea == io_in ? 12'hbce : _GEN_2281; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2283 = 12'h8eb == io_in ? 12'hd80 : _GEN_2282; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2284 = 12'h8ec == io_in ? 12'hd70 : _GEN_2283; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2285 = 12'h8ed == io_in ? 12'h47 : _GEN_2284; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2286 = 12'h8ee == io_in ? 12'hce7 : _GEN_2285; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2287 = 12'h8ef == io_in ? 12'hdca : _GEN_2286; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2288 = 12'h8f0 == io_in ? 12'h9ef : _GEN_2287; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2289 = 12'h8f1 == io_in ? 12'h304 : _GEN_2288; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2290 = 12'h8f2 == io_in ? 12'h116 : _GEN_2289; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2291 = 12'h8f3 == io_in ? 12'h927 : _GEN_2290; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2292 = 12'h8f4 == io_in ? 12'h9f2 : _GEN_2291; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2293 = 12'h8f5 == io_in ? 12'hc84 : _GEN_2292; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2294 = 12'h8f6 == io_in ? 12'h639 : _GEN_2293; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2295 = 12'h8f7 == io_in ? 12'hc3f : _GEN_2294; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2296 = 12'h8f8 == io_in ? 12'he22 : _GEN_2295; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2297 = 12'h8f9 == io_in ? 12'ha08 : _GEN_2296; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2298 = 12'h8fa == io_in ? 12'hf04 : _GEN_2297; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2299 = 12'h8fb == io_in ? 12'he4f : _GEN_2298; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2300 = 12'h8fc == io_in ? 12'hb6e : _GEN_2299; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2301 = 12'h8fd == io_in ? 12'h341 : _GEN_2300; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2302 = 12'h8fe == io_in ? 12'h5b6 : _GEN_2301; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2303 = 12'h8ff == io_in ? 12'hf51 : _GEN_2302; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2304 = 12'h900 == io_in ? 12'h858 : _GEN_2303; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2305 = 12'h901 == io_in ? 12'hc34 : _GEN_2304; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2306 = 12'h902 == io_in ? 12'h8a : _GEN_2305; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2307 = 12'h903 == io_in ? 12'h469 : _GEN_2306; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2308 = 12'h904 == io_in ? 12'h8be : _GEN_2307; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2309 = 12'h905 == io_in ? 12'h272 : _GEN_2308; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2310 = 12'h906 == io_in ? 12'hb26 : _GEN_2309; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2311 = 12'h907 == io_in ? 12'h70d : _GEN_2310; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2312 = 12'h908 == io_in ? 12'h11d : _GEN_2311; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2313 = 12'h909 == io_in ? 12'hd24 : _GEN_2312; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2314 = 12'h90a == io_in ? 12'h464 : _GEN_2313; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2315 = 12'h90b == io_in ? 12'h92e : _GEN_2314; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2316 = 12'h90c == io_in ? 12'ha3e : _GEN_2315; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2317 = 12'h90d == io_in ? 12'h4bd : _GEN_2316; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2318 = 12'h90e == io_in ? 12'hc52 : _GEN_2317; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2319 = 12'h90f == io_in ? 12'hf8e : _GEN_2318; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2320 = 12'h910 == io_in ? 12'h94a : _GEN_2319; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2321 = 12'h911 == io_in ? 12'h5fc : _GEN_2320; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2322 = 12'h912 == io_in ? 12'h3db : _GEN_2321; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2323 = 12'h913 == io_in ? 12'h68c : _GEN_2322; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2324 = 12'h914 == io_in ? 12'h944 : _GEN_2323; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2325 = 12'h915 == io_in ? 12'h78f : _GEN_2324; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2326 = 12'h916 == io_in ? 12'h793 : _GEN_2325; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2327 = 12'h917 == io_in ? 12'h984 : _GEN_2326; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2328 = 12'h918 == io_in ? 12'hf67 : _GEN_2327; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2329 = 12'h919 == io_in ? 12'h791 : _GEN_2328; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2330 = 12'h91a == io_in ? 12'h85f : _GEN_2329; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2331 = 12'h91b == io_in ? 12'h16b : _GEN_2330; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2332 = 12'h91c == io_in ? 12'hcc : _GEN_2331; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2333 = 12'h91d == io_in ? 12'ha62 : _GEN_2332; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2334 = 12'h91e == io_in ? 12'h7ac : _GEN_2333; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2335 = 12'h91f == io_in ? 12'hd36 : _GEN_2334; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2336 = 12'h920 == io_in ? 12'h565 : _GEN_2335; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2337 = 12'h921 == io_in ? 12'h4ec : _GEN_2336; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2338 = 12'h922 == io_in ? 12'he31 : _GEN_2337; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2339 = 12'h923 == io_in ? 12'h285 : _GEN_2338; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2340 = 12'h924 == io_in ? 12'ha10 : _GEN_2339; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2341 = 12'h925 == io_in ? 12'he02 : _GEN_2340; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2342 = 12'h926 == io_in ? 12'hb36 : _GEN_2341; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2343 = 12'h927 == io_in ? 12'h431 : _GEN_2342; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2344 = 12'h928 == io_in ? 12'h411 : _GEN_2343; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2345 = 12'h929 == io_in ? 12'hb42 : _GEN_2344; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2346 = 12'h92a == io_in ? 12'h23b : _GEN_2345; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2347 = 12'h92b == io_in ? 12'hfa6 : _GEN_2346; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2348 = 12'h92c == io_in ? 12'h5ad : _GEN_2347; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2349 = 12'h92d == io_in ? 12'hb43 : _GEN_2348; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2350 = 12'h92e == io_in ? 12'hb16 : _GEN_2349; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2351 = 12'h92f == io_in ? 12'hb5a : _GEN_2350; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2352 = 12'h930 == io_in ? 12'hace : _GEN_2351; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2353 = 12'h931 == io_in ? 12'h782 : _GEN_2352; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2354 = 12'h932 == io_in ? 12'hf64 : _GEN_2353; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2355 = 12'h933 == io_in ? 12'h58d : _GEN_2354; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2356 = 12'h934 == io_in ? 12'h280 : _GEN_2355; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2357 = 12'h935 == io_in ? 12'h219 : _GEN_2356; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2358 = 12'h936 == io_in ? 12'h2f0 : _GEN_2357; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2359 = 12'h937 == io_in ? 12'h11f : _GEN_2358; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2360 = 12'h938 == io_in ? 12'hde4 : _GEN_2359; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2361 = 12'h939 == io_in ? 12'h55a : _GEN_2360; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2362 = 12'h93a == io_in ? 12'hcaf : _GEN_2361; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2363 = 12'h93b == io_in ? 12'hcf : _GEN_2362; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2364 = 12'h93c == io_in ? 12'he38 : _GEN_2363; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2365 = 12'h93d == io_in ? 12'h3ff : _GEN_2364; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2366 = 12'h93e == io_in ? 12'h4af : _GEN_2365; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2367 = 12'h93f == io_in ? 12'h211 : _GEN_2366; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2368 = 12'h940 == io_in ? 12'hbd9 : _GEN_2367; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2369 = 12'h941 == io_in ? 12'hf94 : _GEN_2368; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2370 = 12'h942 == io_in ? 12'h9f : _GEN_2369; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2371 = 12'h943 == io_in ? 12'h700 : _GEN_2370; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2372 = 12'h944 == io_in ? 12'h134 : _GEN_2371; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2373 = 12'h945 == io_in ? 12'h6bd : _GEN_2372; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2374 = 12'h946 == io_in ? 12'h4c8 : _GEN_2373; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2375 = 12'h947 == io_in ? 12'h11c : _GEN_2374; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2376 = 12'h948 == io_in ? 12'hb00 : _GEN_2375; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2377 = 12'h949 == io_in ? 12'h682 : _GEN_2376; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2378 = 12'h94a == io_in ? 12'h842 : _GEN_2377; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2379 = 12'h94b == io_in ? 12'h887 : _GEN_2378; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2380 = 12'h94c == io_in ? 12'h719 : _GEN_2379; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2381 = 12'h94d == io_in ? 12'hfd6 : _GEN_2380; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2382 = 12'h94e == io_in ? 12'hfe7 : _GEN_2381; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2383 = 12'h94f == io_in ? 12'h3c : _GEN_2382; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2384 = 12'h950 == io_in ? 12'hbac : _GEN_2383; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2385 = 12'h951 == io_in ? 12'he18 : _GEN_2384; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2386 = 12'h952 == io_in ? 12'ha5 : _GEN_2385; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2387 = 12'h953 == io_in ? 12'hf66 : _GEN_2386; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2388 = 12'h954 == io_in ? 12'h17 : _GEN_2387; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2389 = 12'h955 == io_in ? 12'h3f2 : _GEN_2388; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2390 = 12'h956 == io_in ? 12'hc65 : _GEN_2389; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2391 = 12'h957 == io_in ? 12'h264 : _GEN_2390; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2392 = 12'h958 == io_in ? 12'h90e : _GEN_2391; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2393 = 12'h959 == io_in ? 12'h32b : _GEN_2392; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2394 = 12'h95a == io_in ? 12'h825 : _GEN_2393; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2395 = 12'h95b == io_in ? 12'hf70 : _GEN_2394; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2396 = 12'h95c == io_in ? 12'hbaf : _GEN_2395; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2397 = 12'h95d == io_in ? 12'h9cd : _GEN_2396; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2398 = 12'h95e == io_in ? 12'h9d7 : _GEN_2397; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2399 = 12'h95f == io_in ? 12'h0 : _GEN_2398; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2400 = 12'h960 == io_in ? 12'h318 : _GEN_2399; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2401 = 12'h961 == io_in ? 12'h55a : _GEN_2400; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2402 = 12'h962 == io_in ? 12'ha84 : _GEN_2401; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2403 = 12'h963 == io_in ? 12'h12e : _GEN_2402; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2404 = 12'h964 == io_in ? 12'hd64 : _GEN_2403; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2405 = 12'h965 == io_in ? 12'hc5d : _GEN_2404; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2406 = 12'h966 == io_in ? 12'hfbf : _GEN_2405; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2407 = 12'h967 == io_in ? 12'h44f : _GEN_2406; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2408 = 12'h968 == io_in ? 12'he5a : _GEN_2407; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2409 = 12'h969 == io_in ? 12'h1bb : _GEN_2408; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2410 = 12'h96a == io_in ? 12'he72 : _GEN_2409; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2411 = 12'h96b == io_in ? 12'h9fe : _GEN_2410; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2412 = 12'h96c == io_in ? 12'h586 : _GEN_2411; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2413 = 12'h96d == io_in ? 12'hce5 : _GEN_2412; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2414 = 12'h96e == io_in ? 12'h94f : _GEN_2413; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2415 = 12'h96f == io_in ? 12'h386 : _GEN_2414; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2416 = 12'h970 == io_in ? 12'hc0b : _GEN_2415; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2417 = 12'h971 == io_in ? 12'h9b0 : _GEN_2416; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2418 = 12'h972 == io_in ? 12'h588 : _GEN_2417; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2419 = 12'h973 == io_in ? 12'h1b5 : _GEN_2418; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2420 = 12'h974 == io_in ? 12'hceb : _GEN_2419; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2421 = 12'h975 == io_in ? 12'h2fb : _GEN_2420; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2422 = 12'h976 == io_in ? 12'h7f6 : _GEN_2421; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2423 = 12'h977 == io_in ? 12'hf86 : _GEN_2422; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2424 = 12'h978 == io_in ? 12'h42a : _GEN_2423; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2425 = 12'h979 == io_in ? 12'hc9 : _GEN_2424; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2426 = 12'h97a == io_in ? 12'h90 : _GEN_2425; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2427 = 12'h97b == io_in ? 12'h856 : _GEN_2426; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2428 = 12'h97c == io_in ? 12'h13a : _GEN_2427; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2429 = 12'h97d == io_in ? 12'he85 : _GEN_2428; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2430 = 12'h97e == io_in ? 12'h58 : _GEN_2429; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2431 = 12'h97f == io_in ? 12'h38f : _GEN_2430; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2432 = 12'h980 == io_in ? 12'h5d5 : _GEN_2431; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2433 = 12'h981 == io_in ? 12'hcc2 : _GEN_2432; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2434 = 12'h982 == io_in ? 12'h146 : _GEN_2433; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2435 = 12'h983 == io_in ? 12'h527 : _GEN_2434; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2436 = 12'h984 == io_in ? 12'h8ea : _GEN_2435; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2437 = 12'h985 == io_in ? 12'hdf8 : _GEN_2436; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2438 = 12'h986 == io_in ? 12'hdfc : _GEN_2437; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2439 = 12'h987 == io_in ? 12'he59 : _GEN_2438; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2440 = 12'h988 == io_in ? 12'he94 : _GEN_2439; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2441 = 12'h989 == io_in ? 12'h370 : _GEN_2440; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2442 = 12'h98a == io_in ? 12'h90 : _GEN_2441; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2443 = 12'h98b == io_in ? 12'h3d0 : _GEN_2442; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2444 = 12'h98c == io_in ? 12'ha1a : _GEN_2443; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2445 = 12'h98d == io_in ? 12'h219 : _GEN_2444; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2446 = 12'h98e == io_in ? 12'h10b : _GEN_2445; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2447 = 12'h98f == io_in ? 12'hd6b : _GEN_2446; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2448 = 12'h990 == io_in ? 12'h8ac : _GEN_2447; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2449 = 12'h991 == io_in ? 12'h363 : _GEN_2448; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2450 = 12'h992 == io_in ? 12'h480 : _GEN_2449; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2451 = 12'h993 == io_in ? 12'h3c4 : _GEN_2450; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2452 = 12'h994 == io_in ? 12'hdc4 : _GEN_2451; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2453 = 12'h995 == io_in ? 12'h7dd : _GEN_2452; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2454 = 12'h996 == io_in ? 12'hf07 : _GEN_2453; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2455 = 12'h997 == io_in ? 12'h4bb : _GEN_2454; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2456 = 12'h998 == io_in ? 12'h22e : _GEN_2455; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2457 = 12'h999 == io_in ? 12'h5c4 : _GEN_2456; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2458 = 12'h99a == io_in ? 12'hc4f : _GEN_2457; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2459 = 12'h99b == io_in ? 12'h2aa : _GEN_2458; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2460 = 12'h99c == io_in ? 12'h1d1 : _GEN_2459; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2461 = 12'h99d == io_in ? 12'h8fb : _GEN_2460; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2462 = 12'h99e == io_in ? 12'h384 : _GEN_2461; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2463 = 12'h99f == io_in ? 12'h1e3 : _GEN_2462; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2464 = 12'h9a0 == io_in ? 12'h29f : _GEN_2463; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2465 = 12'h9a1 == io_in ? 12'ha26 : _GEN_2464; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2466 = 12'h9a2 == io_in ? 12'h9bf : _GEN_2465; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2467 = 12'h9a3 == io_in ? 12'h31e : _GEN_2466; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2468 = 12'h9a4 == io_in ? 12'hff8 : _GEN_2467; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2469 = 12'h9a5 == io_in ? 12'h3fd : _GEN_2468; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2470 = 12'h9a6 == io_in ? 12'h77 : _GEN_2469; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2471 = 12'h9a7 == io_in ? 12'hb83 : _GEN_2470; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2472 = 12'h9a8 == io_in ? 12'hbeb : _GEN_2471; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2473 = 12'h9a9 == io_in ? 12'hf7a : _GEN_2472; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2474 = 12'h9aa == io_in ? 12'h73f : _GEN_2473; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2475 = 12'h9ab == io_in ? 12'he75 : _GEN_2474; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2476 = 12'h9ac == io_in ? 12'hd6c : _GEN_2475; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2477 = 12'h9ad == io_in ? 12'h5b9 : _GEN_2476; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2478 = 12'h9ae == io_in ? 12'hebd : _GEN_2477; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2479 = 12'h9af == io_in ? 12'haac : _GEN_2478; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2480 = 12'h9b0 == io_in ? 12'hc65 : _GEN_2479; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2481 = 12'h9b1 == io_in ? 12'hab : _GEN_2480; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2482 = 12'h9b2 == io_in ? 12'h870 : _GEN_2481; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2483 = 12'h9b3 == io_in ? 12'h1e6 : _GEN_2482; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2484 = 12'h9b4 == io_in ? 12'hf8c : _GEN_2483; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2485 = 12'h9b5 == io_in ? 12'hf50 : _GEN_2484; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2486 = 12'h9b6 == io_in ? 12'hf1f : _GEN_2485; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2487 = 12'h9b7 == io_in ? 12'h66d : _GEN_2486; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2488 = 12'h9b8 == io_in ? 12'h366 : _GEN_2487; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2489 = 12'h9b9 == io_in ? 12'hee2 : _GEN_2488; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2490 = 12'h9ba == io_in ? 12'h787 : _GEN_2489; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2491 = 12'h9bb == io_in ? 12'hddc : _GEN_2490; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2492 = 12'h9bc == io_in ? 12'h50f : _GEN_2491; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2493 = 12'h9bd == io_in ? 12'hdc5 : _GEN_2492; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2494 = 12'h9be == io_in ? 12'ha29 : _GEN_2493; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2495 = 12'h9bf == io_in ? 12'hfe8 : _GEN_2494; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2496 = 12'h9c0 == io_in ? 12'h842 : _GEN_2495; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2497 = 12'h9c1 == io_in ? 12'h7b9 : _GEN_2496; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2498 = 12'h9c2 == io_in ? 12'hd4c : _GEN_2497; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2499 = 12'h9c3 == io_in ? 12'h8c7 : _GEN_2498; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2500 = 12'h9c4 == io_in ? 12'h55 : _GEN_2499; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2501 = 12'h9c5 == io_in ? 12'habd : _GEN_2500; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2502 = 12'h9c6 == io_in ? 12'h9aa : _GEN_2501; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2503 = 12'h9c7 == io_in ? 12'h87 : _GEN_2502; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2504 = 12'h9c8 == io_in ? 12'h3fb : _GEN_2503; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2505 = 12'h9c9 == io_in ? 12'ha2b : _GEN_2504; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2506 = 12'h9ca == io_in ? 12'h368 : _GEN_2505; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2507 = 12'h9cb == io_in ? 12'h642 : _GEN_2506; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2508 = 12'h9cc == io_in ? 12'h79f : _GEN_2507; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2509 = 12'h9cd == io_in ? 12'h89c : _GEN_2508; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2510 = 12'h9ce == io_in ? 12'h1e3 : _GEN_2509; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2511 = 12'h9cf == io_in ? 12'hb52 : _GEN_2510; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2512 = 12'h9d0 == io_in ? 12'h163 : _GEN_2511; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2513 = 12'h9d1 == io_in ? 12'h23c : _GEN_2512; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2514 = 12'h9d2 == io_in ? 12'h8e6 : _GEN_2513; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2515 = 12'h9d3 == io_in ? 12'h6ef : _GEN_2514; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2516 = 12'h9d4 == io_in ? 12'h261 : _GEN_2515; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2517 = 12'h9d5 == io_in ? 12'hfe7 : _GEN_2516; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2518 = 12'h9d6 == io_in ? 12'h9f8 : _GEN_2517; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2519 = 12'h9d7 == io_in ? 12'he79 : _GEN_2518; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2520 = 12'h9d8 == io_in ? 12'hcf3 : _GEN_2519; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2521 = 12'h9d9 == io_in ? 12'h914 : _GEN_2520; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2522 = 12'h9da == io_in ? 12'hfae : _GEN_2521; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2523 = 12'h9db == io_in ? 12'hdd7 : _GEN_2522; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2524 = 12'h9dc == io_in ? 12'h7bc : _GEN_2523; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2525 = 12'h9dd == io_in ? 12'hf78 : _GEN_2524; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2526 = 12'h9de == io_in ? 12'hb2e : _GEN_2525; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2527 = 12'h9df == io_in ? 12'ha99 : _GEN_2526; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2528 = 12'h9e0 == io_in ? 12'h5f2 : _GEN_2527; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2529 = 12'h9e1 == io_in ? 12'hd29 : _GEN_2528; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2530 = 12'h9e2 == io_in ? 12'hf2a : _GEN_2529; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2531 = 12'h9e3 == io_in ? 12'h4d0 : _GEN_2530; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2532 = 12'h9e4 == io_in ? 12'h9d0 : _GEN_2531; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2533 = 12'h9e5 == io_in ? 12'h58b : _GEN_2532; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2534 = 12'h9e6 == io_in ? 12'h546 : _GEN_2533; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2535 = 12'h9e7 == io_in ? 12'ha5a : _GEN_2534; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2536 = 12'h9e8 == io_in ? 12'hd1b : _GEN_2535; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2537 = 12'h9e9 == io_in ? 12'hd11 : _GEN_2536; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2538 = 12'h9ea == io_in ? 12'h3eb : _GEN_2537; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2539 = 12'h9eb == io_in ? 12'haa7 : _GEN_2538; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2540 = 12'h9ec == io_in ? 12'hb51 : _GEN_2539; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2541 = 12'h9ed == io_in ? 12'h4a2 : _GEN_2540; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2542 = 12'h9ee == io_in ? 12'hb2c : _GEN_2541; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2543 = 12'h9ef == io_in ? 12'h680 : _GEN_2542; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2544 = 12'h9f0 == io_in ? 12'ha42 : _GEN_2543; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2545 = 12'h9f1 == io_in ? 12'h666 : _GEN_2544; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2546 = 12'h9f2 == io_in ? 12'h69e : _GEN_2545; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2547 = 12'h9f3 == io_in ? 12'hba8 : _GEN_2546; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2548 = 12'h9f4 == io_in ? 12'h976 : _GEN_2547; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2549 = 12'h9f5 == io_in ? 12'hc7e : _GEN_2548; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2550 = 12'h9f6 == io_in ? 12'hee1 : _GEN_2549; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2551 = 12'h9f7 == io_in ? 12'h83 : _GEN_2550; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2552 = 12'h9f8 == io_in ? 12'h212 : _GEN_2551; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2553 = 12'h9f9 == io_in ? 12'h1fa : _GEN_2552; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2554 = 12'h9fa == io_in ? 12'hd6d : _GEN_2553; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2555 = 12'h9fb == io_in ? 12'hf41 : _GEN_2554; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2556 = 12'h9fc == io_in ? 12'hb1a : _GEN_2555; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2557 = 12'h9fd == io_in ? 12'hd68 : _GEN_2556; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2558 = 12'h9fe == io_in ? 12'h58d : _GEN_2557; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2559 = 12'h9ff == io_in ? 12'h856 : _GEN_2558; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2560 = 12'ha00 == io_in ? 12'h74e : _GEN_2559; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2561 = 12'ha01 == io_in ? 12'hec0 : _GEN_2560; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2562 = 12'ha02 == io_in ? 12'ha2d : _GEN_2561; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2563 = 12'ha03 == io_in ? 12'h465 : _GEN_2562; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2564 = 12'ha04 == io_in ? 12'h78c : _GEN_2563; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2565 = 12'ha05 == io_in ? 12'h265 : _GEN_2564; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2566 = 12'ha06 == io_in ? 12'hd44 : _GEN_2565; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2567 = 12'ha07 == io_in ? 12'h907 : _GEN_2566; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2568 = 12'ha08 == io_in ? 12'h796 : _GEN_2567; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2569 = 12'ha09 == io_in ? 12'h547 : _GEN_2568; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2570 = 12'ha0a == io_in ? 12'hda1 : _GEN_2569; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2571 = 12'ha0b == io_in ? 12'h977 : _GEN_2570; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2572 = 12'ha0c == io_in ? 12'h354 : _GEN_2571; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2573 = 12'ha0d == io_in ? 12'hdcd : _GEN_2572; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2574 = 12'ha0e == io_in ? 12'hd0f : _GEN_2573; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2575 = 12'ha0f == io_in ? 12'hb4e : _GEN_2574; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2576 = 12'ha10 == io_in ? 12'haf6 : _GEN_2575; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2577 = 12'ha11 == io_in ? 12'h700 : _GEN_2576; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2578 = 12'ha12 == io_in ? 12'h45e : _GEN_2577; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2579 = 12'ha13 == io_in ? 12'h467 : _GEN_2578; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2580 = 12'ha14 == io_in ? 12'h7c5 : _GEN_2579; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2581 = 12'ha15 == io_in ? 12'hb26 : _GEN_2580; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2582 = 12'ha16 == io_in ? 12'h56f : _GEN_2581; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2583 = 12'ha17 == io_in ? 12'hd54 : _GEN_2582; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2584 = 12'ha18 == io_in ? 12'h739 : _GEN_2583; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2585 = 12'ha19 == io_in ? 12'h5fe : _GEN_2584; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2586 = 12'ha1a == io_in ? 12'h4c5 : _GEN_2585; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2587 = 12'ha1b == io_in ? 12'hbd1 : _GEN_2586; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2588 = 12'ha1c == io_in ? 12'hb0e : _GEN_2587; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2589 = 12'ha1d == io_in ? 12'h909 : _GEN_2588; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2590 = 12'ha1e == io_in ? 12'h398 : _GEN_2589; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2591 = 12'ha1f == io_in ? 12'hb4a : _GEN_2590; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2592 = 12'ha20 == io_in ? 12'h42c : _GEN_2591; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2593 = 12'ha21 == io_in ? 12'hc27 : _GEN_2592; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2594 = 12'ha22 == io_in ? 12'heb7 : _GEN_2593; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2595 = 12'ha23 == io_in ? 12'h2cb : _GEN_2594; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2596 = 12'ha24 == io_in ? 12'ha18 : _GEN_2595; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2597 = 12'ha25 == io_in ? 12'h633 : _GEN_2596; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2598 = 12'ha26 == io_in ? 12'h439 : _GEN_2597; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2599 = 12'ha27 == io_in ? 12'hd92 : _GEN_2598; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2600 = 12'ha28 == io_in ? 12'hca9 : _GEN_2599; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2601 = 12'ha29 == io_in ? 12'h34d : _GEN_2600; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2602 = 12'ha2a == io_in ? 12'hdb2 : _GEN_2601; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2603 = 12'ha2b == io_in ? 12'he44 : _GEN_2602; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2604 = 12'ha2c == io_in ? 12'hb3e : _GEN_2603; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2605 = 12'ha2d == io_in ? 12'hddb : _GEN_2604; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2606 = 12'ha2e == io_in ? 12'hbbd : _GEN_2605; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2607 = 12'ha2f == io_in ? 12'h6b3 : _GEN_2606; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2608 = 12'ha30 == io_in ? 12'h97e : _GEN_2607; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2609 = 12'ha31 == io_in ? 12'haf2 : _GEN_2608; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2610 = 12'ha32 == io_in ? 12'h41d : _GEN_2609; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2611 = 12'ha33 == io_in ? 12'h4aa : _GEN_2610; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2612 = 12'ha34 == io_in ? 12'h18d : _GEN_2611; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2613 = 12'ha35 == io_in ? 12'h8af : _GEN_2612; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2614 = 12'ha36 == io_in ? 12'h181 : _GEN_2613; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2615 = 12'ha37 == io_in ? 12'hd4d : _GEN_2614; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2616 = 12'ha38 == io_in ? 12'h701 : _GEN_2615; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2617 = 12'ha39 == io_in ? 12'h3f4 : _GEN_2616; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2618 = 12'ha3a == io_in ? 12'h38f : _GEN_2617; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2619 = 12'ha3b == io_in ? 12'h6b1 : _GEN_2618; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2620 = 12'ha3c == io_in ? 12'h315 : _GEN_2619; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2621 = 12'ha3d == io_in ? 12'h9d0 : _GEN_2620; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2622 = 12'ha3e == io_in ? 12'h18d : _GEN_2621; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2623 = 12'ha3f == io_in ? 12'hcdb : _GEN_2622; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2624 = 12'ha40 == io_in ? 12'hc37 : _GEN_2623; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2625 = 12'ha41 == io_in ? 12'h6a9 : _GEN_2624; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2626 = 12'ha42 == io_in ? 12'h90e : _GEN_2625; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2627 = 12'ha43 == io_in ? 12'h304 : _GEN_2626; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2628 = 12'ha44 == io_in ? 12'ha59 : _GEN_2627; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2629 = 12'ha45 == io_in ? 12'h98f : _GEN_2628; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2630 = 12'ha46 == io_in ? 12'hd00 : _GEN_2629; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2631 = 12'ha47 == io_in ? 12'h2f9 : _GEN_2630; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2632 = 12'ha48 == io_in ? 12'h356 : _GEN_2631; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2633 = 12'ha49 == io_in ? 12'h47b : _GEN_2632; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2634 = 12'ha4a == io_in ? 12'he3a : _GEN_2633; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2635 = 12'ha4b == io_in ? 12'hdcc : _GEN_2634; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2636 = 12'ha4c == io_in ? 12'hac3 : _GEN_2635; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2637 = 12'ha4d == io_in ? 12'h278 : _GEN_2636; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2638 = 12'ha4e == io_in ? 12'h45d : _GEN_2637; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2639 = 12'ha4f == io_in ? 12'h688 : _GEN_2638; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2640 = 12'ha50 == io_in ? 12'he6f : _GEN_2639; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2641 = 12'ha51 == io_in ? 12'h346 : _GEN_2640; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2642 = 12'ha52 == io_in ? 12'h77 : _GEN_2641; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2643 = 12'ha53 == io_in ? 12'hc6 : _GEN_2642; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2644 = 12'ha54 == io_in ? 12'haa4 : _GEN_2643; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2645 = 12'ha55 == io_in ? 12'hb6 : _GEN_2644; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2646 = 12'ha56 == io_in ? 12'h88f : _GEN_2645; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2647 = 12'ha57 == io_in ? 12'h9e9 : _GEN_2646; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2648 = 12'ha58 == io_in ? 12'he1 : _GEN_2647; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2649 = 12'ha59 == io_in ? 12'he56 : _GEN_2648; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2650 = 12'ha5a == io_in ? 12'h644 : _GEN_2649; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2651 = 12'ha5b == io_in ? 12'h8f0 : _GEN_2650; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2652 = 12'ha5c == io_in ? 12'ha08 : _GEN_2651; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2653 = 12'ha5d == io_in ? 12'h7b0 : _GEN_2652; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2654 = 12'ha5e == io_in ? 12'hf7f : _GEN_2653; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2655 = 12'ha5f == io_in ? 12'ha35 : _GEN_2654; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2656 = 12'ha60 == io_in ? 12'h660 : _GEN_2655; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2657 = 12'ha61 == io_in ? 12'h713 : _GEN_2656; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2658 = 12'ha62 == io_in ? 12'h7fa : _GEN_2657; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2659 = 12'ha63 == io_in ? 12'hb8a : _GEN_2658; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2660 = 12'ha64 == io_in ? 12'hd3f : _GEN_2659; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2661 = 12'ha65 == io_in ? 12'he26 : _GEN_2660; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2662 = 12'ha66 == io_in ? 12'h7b6 : _GEN_2661; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2663 = 12'ha67 == io_in ? 12'ha39 : _GEN_2662; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2664 = 12'ha68 == io_in ? 12'h30b : _GEN_2663; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2665 = 12'ha69 == io_in ? 12'hdfb : _GEN_2664; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2666 = 12'ha6a == io_in ? 12'h539 : _GEN_2665; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2667 = 12'ha6b == io_in ? 12'h572 : _GEN_2666; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2668 = 12'ha6c == io_in ? 12'hbe4 : _GEN_2667; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2669 = 12'ha6d == io_in ? 12'h5ff : _GEN_2668; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2670 = 12'ha6e == io_in ? 12'h399 : _GEN_2669; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2671 = 12'ha6f == io_in ? 12'h192 : _GEN_2670; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2672 = 12'ha70 == io_in ? 12'hd45 : _GEN_2671; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2673 = 12'ha71 == io_in ? 12'hbc3 : _GEN_2672; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2674 = 12'ha72 == io_in ? 12'ha79 : _GEN_2673; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2675 = 12'ha73 == io_in ? 12'h5a7 : _GEN_2674; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2676 = 12'ha74 == io_in ? 12'h999 : _GEN_2675; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2677 = 12'ha75 == io_in ? 12'h251 : _GEN_2676; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2678 = 12'ha76 == io_in ? 12'h4d : _GEN_2677; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2679 = 12'ha77 == io_in ? 12'he4c : _GEN_2678; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2680 = 12'ha78 == io_in ? 12'h9b7 : _GEN_2679; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2681 = 12'ha79 == io_in ? 12'h204 : _GEN_2680; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2682 = 12'ha7a == io_in ? 12'hb1c : _GEN_2681; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2683 = 12'ha7b == io_in ? 12'h607 : _GEN_2682; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2684 = 12'ha7c == io_in ? 12'hcad : _GEN_2683; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2685 = 12'ha7d == io_in ? 12'h420 : _GEN_2684; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2686 = 12'ha7e == io_in ? 12'h688 : _GEN_2685; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2687 = 12'ha7f == io_in ? 12'h9dd : _GEN_2686; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2688 = 12'ha80 == io_in ? 12'hc1a : _GEN_2687; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2689 = 12'ha81 == io_in ? 12'hb19 : _GEN_2688; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2690 = 12'ha82 == io_in ? 12'hbb0 : _GEN_2689; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2691 = 12'ha83 == io_in ? 12'hc10 : _GEN_2690; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2692 = 12'ha84 == io_in ? 12'h50 : _GEN_2691; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2693 = 12'ha85 == io_in ? 12'h4a1 : _GEN_2692; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2694 = 12'ha86 == io_in ? 12'hc04 : _GEN_2693; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2695 = 12'ha87 == io_in ? 12'h165 : _GEN_2694; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2696 = 12'ha88 == io_in ? 12'hc0f : _GEN_2695; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2697 = 12'ha89 == io_in ? 12'h15d : _GEN_2696; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2698 = 12'ha8a == io_in ? 12'h5d8 : _GEN_2697; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2699 = 12'ha8b == io_in ? 12'h6c9 : _GEN_2698; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2700 = 12'ha8c == io_in ? 12'h3e9 : _GEN_2699; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2701 = 12'ha8d == io_in ? 12'hac8 : _GEN_2700; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2702 = 12'ha8e == io_in ? 12'h37e : _GEN_2701; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2703 = 12'ha8f == io_in ? 12'hc9e : _GEN_2702; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2704 = 12'ha90 == io_in ? 12'hc8e : _GEN_2703; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2705 = 12'ha91 == io_in ? 12'h72a : _GEN_2704; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2706 = 12'ha92 == io_in ? 12'h3b4 : _GEN_2705; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2707 = 12'ha93 == io_in ? 12'hea0 : _GEN_2706; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2708 = 12'ha94 == io_in ? 12'h7a0 : _GEN_2707; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2709 = 12'ha95 == io_in ? 12'h93c : _GEN_2708; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2710 = 12'ha96 == io_in ? 12'he9d : _GEN_2709; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2711 = 12'ha97 == io_in ? 12'h6e6 : _GEN_2710; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2712 = 12'ha98 == io_in ? 12'h626 : _GEN_2711; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2713 = 12'ha99 == io_in ? 12'haa1 : _GEN_2712; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2714 = 12'ha9a == io_in ? 12'hb78 : _GEN_2713; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2715 = 12'ha9b == io_in ? 12'h6b : _GEN_2714; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2716 = 12'ha9c == io_in ? 12'hf23 : _GEN_2715; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2717 = 12'ha9d == io_in ? 12'h9b2 : _GEN_2716; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2718 = 12'ha9e == io_in ? 12'h951 : _GEN_2717; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2719 = 12'ha9f == io_in ? 12'h255 : _GEN_2718; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2720 = 12'haa0 == io_in ? 12'h86d : _GEN_2719; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2721 = 12'haa1 == io_in ? 12'h254 : _GEN_2720; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2722 = 12'haa2 == io_in ? 12'h51b : _GEN_2721; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2723 = 12'haa3 == io_in ? 12'h55e : _GEN_2722; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2724 = 12'haa4 == io_in ? 12'h703 : _GEN_2723; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2725 = 12'haa5 == io_in ? 12'hb20 : _GEN_2724; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2726 = 12'haa6 == io_in ? 12'h8b4 : _GEN_2725; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2727 = 12'haa7 == io_in ? 12'hdd4 : _GEN_2726; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2728 = 12'haa8 == io_in ? 12'hdc8 : _GEN_2727; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2729 = 12'haa9 == io_in ? 12'h2ad : _GEN_2728; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2730 = 12'haaa == io_in ? 12'hbfe : _GEN_2729; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2731 = 12'haab == io_in ? 12'h730 : _GEN_2730; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2732 = 12'haac == io_in ? 12'h730 : _GEN_2731; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2733 = 12'haad == io_in ? 12'h10a : _GEN_2732; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2734 = 12'haae == io_in ? 12'h8a6 : _GEN_2733; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2735 = 12'haaf == io_in ? 12'h4af : _GEN_2734; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2736 = 12'hab0 == io_in ? 12'h5e0 : _GEN_2735; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2737 = 12'hab1 == io_in ? 12'heef : _GEN_2736; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2738 = 12'hab2 == io_in ? 12'hcac : _GEN_2737; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2739 = 12'hab3 == io_in ? 12'h149 : _GEN_2738; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2740 = 12'hab4 == io_in ? 12'h55a : _GEN_2739; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2741 = 12'hab5 == io_in ? 12'h3a0 : _GEN_2740; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2742 = 12'hab6 == io_in ? 12'h2cf : _GEN_2741; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2743 = 12'hab7 == io_in ? 12'h821 : _GEN_2742; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2744 = 12'hab8 == io_in ? 12'h6bc : _GEN_2743; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2745 = 12'hab9 == io_in ? 12'hc73 : _GEN_2744; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2746 = 12'haba == io_in ? 12'h39e : _GEN_2745; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2747 = 12'habb == io_in ? 12'h631 : _GEN_2746; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2748 = 12'habc == io_in ? 12'hd0f : _GEN_2747; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2749 = 12'habd == io_in ? 12'ha3e : _GEN_2748; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2750 = 12'habe == io_in ? 12'h7e7 : _GEN_2749; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2751 = 12'habf == io_in ? 12'h9d1 : _GEN_2750; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2752 = 12'hac0 == io_in ? 12'h2cd : _GEN_2751; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2753 = 12'hac1 == io_in ? 12'h2ca : _GEN_2752; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2754 = 12'hac2 == io_in ? 12'hd61 : _GEN_2753; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2755 = 12'hac3 == io_in ? 12'hb39 : _GEN_2754; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2756 = 12'hac4 == io_in ? 12'he3 : _GEN_2755; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2757 = 12'hac5 == io_in ? 12'hc4c : _GEN_2756; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2758 = 12'hac6 == io_in ? 12'ha0 : _GEN_2757; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2759 = 12'hac7 == io_in ? 12'h156 : _GEN_2758; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2760 = 12'hac8 == io_in ? 12'h2ce : _GEN_2759; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2761 = 12'hac9 == io_in ? 12'h829 : _GEN_2760; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2762 = 12'haca == io_in ? 12'ha33 : _GEN_2761; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2763 = 12'hacb == io_in ? 12'hb80 : _GEN_2762; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2764 = 12'hacc == io_in ? 12'hfca : _GEN_2763; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2765 = 12'hacd == io_in ? 12'hf4c : _GEN_2764; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2766 = 12'hace == io_in ? 12'h6ba : _GEN_2765; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2767 = 12'hacf == io_in ? 12'h63e : _GEN_2766; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2768 = 12'had0 == io_in ? 12'h59e : _GEN_2767; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2769 = 12'had1 == io_in ? 12'he8f : _GEN_2768; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2770 = 12'had2 == io_in ? 12'hf86 : _GEN_2769; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2771 = 12'had3 == io_in ? 12'h76d : _GEN_2770; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2772 = 12'had4 == io_in ? 12'hc5d : _GEN_2771; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2773 = 12'had5 == io_in ? 12'hc68 : _GEN_2772; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2774 = 12'had6 == io_in ? 12'h34 : _GEN_2773; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2775 = 12'had7 == io_in ? 12'h427 : _GEN_2774; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2776 = 12'had8 == io_in ? 12'hdf1 : _GEN_2775; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2777 = 12'had9 == io_in ? 12'hbdc : _GEN_2776; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2778 = 12'hada == io_in ? 12'hc2 : _GEN_2777; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2779 = 12'hadb == io_in ? 12'hdc1 : _GEN_2778; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2780 = 12'hadc == io_in ? 12'ha6 : _GEN_2779; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2781 = 12'hadd == io_in ? 12'h398 : _GEN_2780; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2782 = 12'hade == io_in ? 12'hee0 : _GEN_2781; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2783 = 12'hadf == io_in ? 12'h6ff : _GEN_2782; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2784 = 12'hae0 == io_in ? 12'hdd1 : _GEN_2783; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2785 = 12'hae1 == io_in ? 12'hd09 : _GEN_2784; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2786 = 12'hae2 == io_in ? 12'hdcb : _GEN_2785; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2787 = 12'hae3 == io_in ? 12'h853 : _GEN_2786; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2788 = 12'hae4 == io_in ? 12'h8d : _GEN_2787; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2789 = 12'hae5 == io_in ? 12'h6eb : _GEN_2788; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2790 = 12'hae6 == io_in ? 12'hce9 : _GEN_2789; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2791 = 12'hae7 == io_in ? 12'h282 : _GEN_2790; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2792 = 12'hae8 == io_in ? 12'hac9 : _GEN_2791; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2793 = 12'hae9 == io_in ? 12'hb7b : _GEN_2792; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2794 = 12'haea == io_in ? 12'h1d1 : _GEN_2793; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2795 = 12'haeb == io_in ? 12'h7c0 : _GEN_2794; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2796 = 12'haec == io_in ? 12'hee5 : _GEN_2795; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2797 = 12'haed == io_in ? 12'h561 : _GEN_2796; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2798 = 12'haee == io_in ? 12'h43a : _GEN_2797; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2799 = 12'haef == io_in ? 12'h983 : _GEN_2798; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2800 = 12'haf0 == io_in ? 12'h290 : _GEN_2799; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2801 = 12'haf1 == io_in ? 12'h274 : _GEN_2800; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2802 = 12'haf2 == io_in ? 12'hf19 : _GEN_2801; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2803 = 12'haf3 == io_in ? 12'hf0d : _GEN_2802; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2804 = 12'haf4 == io_in ? 12'h59b : _GEN_2803; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2805 = 12'haf5 == io_in ? 12'h224 : _GEN_2804; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2806 = 12'haf6 == io_in ? 12'h1ff : _GEN_2805; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2807 = 12'haf7 == io_in ? 12'h7af : _GEN_2806; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2808 = 12'haf8 == io_in ? 12'h7ed : _GEN_2807; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2809 = 12'haf9 == io_in ? 12'ha62 : _GEN_2808; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2810 = 12'hafa == io_in ? 12'hd68 : _GEN_2809; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2811 = 12'hafb == io_in ? 12'ha97 : _GEN_2810; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2812 = 12'hafc == io_in ? 12'h87e : _GEN_2811; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2813 = 12'hafd == io_in ? 12'h2d8 : _GEN_2812; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2814 = 12'hafe == io_in ? 12'h9d1 : _GEN_2813; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2815 = 12'haff == io_in ? 12'hadb : _GEN_2814; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2816 = 12'hb00 == io_in ? 12'h1ad : _GEN_2815; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2817 = 12'hb01 == io_in ? 12'h7d1 : _GEN_2816; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2818 = 12'hb02 == io_in ? 12'hff2 : _GEN_2817; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2819 = 12'hb03 == io_in ? 12'hc5c : _GEN_2818; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2820 = 12'hb04 == io_in ? 12'hb74 : _GEN_2819; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2821 = 12'hb05 == io_in ? 12'h613 : _GEN_2820; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2822 = 12'hb06 == io_in ? 12'hc81 : _GEN_2821; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2823 = 12'hb07 == io_in ? 12'h9 : _GEN_2822; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2824 = 12'hb08 == io_in ? 12'ha2b : _GEN_2823; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2825 = 12'hb09 == io_in ? 12'h487 : _GEN_2824; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2826 = 12'hb0a == io_in ? 12'hd8c : _GEN_2825; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2827 = 12'hb0b == io_in ? 12'haf7 : _GEN_2826; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2828 = 12'hb0c == io_in ? 12'h108 : _GEN_2827; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2829 = 12'hb0d == io_in ? 12'h1fc : _GEN_2828; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2830 = 12'hb0e == io_in ? 12'h5a2 : _GEN_2829; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2831 = 12'hb0f == io_in ? 12'hbd4 : _GEN_2830; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2832 = 12'hb10 == io_in ? 12'h549 : _GEN_2831; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2833 = 12'hb11 == io_in ? 12'h262 : _GEN_2832; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2834 = 12'hb12 == io_in ? 12'h23d : _GEN_2833; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2835 = 12'hb13 == io_in ? 12'h86a : _GEN_2834; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2836 = 12'hb14 == io_in ? 12'hc92 : _GEN_2835; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2837 = 12'hb15 == io_in ? 12'h27e : _GEN_2836; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2838 = 12'hb16 == io_in ? 12'h76 : _GEN_2837; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2839 = 12'hb17 == io_in ? 12'h5e1 : _GEN_2838; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2840 = 12'hb18 == io_in ? 12'hc2a : _GEN_2839; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2841 = 12'hb19 == io_in ? 12'h140 : _GEN_2840; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2842 = 12'hb1a == io_in ? 12'h408 : _GEN_2841; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2843 = 12'hb1b == io_in ? 12'h21a : _GEN_2842; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2844 = 12'hb1c == io_in ? 12'h436 : _GEN_2843; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2845 = 12'hb1d == io_in ? 12'he35 : _GEN_2844; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2846 = 12'hb1e == io_in ? 12'h114 : _GEN_2845; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2847 = 12'hb1f == io_in ? 12'hb8f : _GEN_2846; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2848 = 12'hb20 == io_in ? 12'ha7f : _GEN_2847; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2849 = 12'hb21 == io_in ? 12'hb4d : _GEN_2848; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2850 = 12'hb22 == io_in ? 12'he3a : _GEN_2849; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2851 = 12'hb23 == io_in ? 12'hc12 : _GEN_2850; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2852 = 12'hb24 == io_in ? 12'ha7d : _GEN_2851; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2853 = 12'hb25 == io_in ? 12'h1e1 : _GEN_2852; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2854 = 12'hb26 == io_in ? 12'h904 : _GEN_2853; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2855 = 12'hb27 == io_in ? 12'h723 : _GEN_2854; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2856 = 12'hb28 == io_in ? 12'h7ad : _GEN_2855; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2857 = 12'hb29 == io_in ? 12'h5cb : _GEN_2856; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2858 = 12'hb2a == io_in ? 12'h643 : _GEN_2857; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2859 = 12'hb2b == io_in ? 12'hf03 : _GEN_2858; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2860 = 12'hb2c == io_in ? 12'hd26 : _GEN_2859; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2861 = 12'hb2d == io_in ? 12'h2d0 : _GEN_2860; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2862 = 12'hb2e == io_in ? 12'h7d0 : _GEN_2861; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2863 = 12'hb2f == io_in ? 12'he12 : _GEN_2862; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2864 = 12'hb30 == io_in ? 12'h75d : _GEN_2863; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2865 = 12'hb31 == io_in ? 12'hf7e : _GEN_2864; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2866 = 12'hb32 == io_in ? 12'h37a : _GEN_2865; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2867 = 12'hb33 == io_in ? 12'ha29 : _GEN_2866; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2868 = 12'hb34 == io_in ? 12'h749 : _GEN_2867; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2869 = 12'hb35 == io_in ? 12'h23b : _GEN_2868; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2870 = 12'hb36 == io_in ? 12'hf77 : _GEN_2869; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2871 = 12'hb37 == io_in ? 12'hb43 : _GEN_2870; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2872 = 12'hb38 == io_in ? 12'hd4 : _GEN_2871; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2873 = 12'hb39 == io_in ? 12'h191 : _GEN_2872; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2874 = 12'hb3a == io_in ? 12'hf : _GEN_2873; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2875 = 12'hb3b == io_in ? 12'h87c : _GEN_2874; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2876 = 12'hb3c == io_in ? 12'hfe8 : _GEN_2875; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2877 = 12'hb3d == io_in ? 12'hd67 : _GEN_2876; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2878 = 12'hb3e == io_in ? 12'hadd : _GEN_2877; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2879 = 12'hb3f == io_in ? 12'h872 : _GEN_2878; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2880 = 12'hb40 == io_in ? 12'h275 : _GEN_2879; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2881 = 12'hb41 == io_in ? 12'h3df : _GEN_2880; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2882 = 12'hb42 == io_in ? 12'hcaa : _GEN_2881; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2883 = 12'hb43 == io_in ? 12'hb69 : _GEN_2882; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2884 = 12'hb44 == io_in ? 12'h368 : _GEN_2883; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2885 = 12'hb45 == io_in ? 12'hca : _GEN_2884; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2886 = 12'hb46 == io_in ? 12'h8e3 : _GEN_2885; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2887 = 12'hb47 == io_in ? 12'h507 : _GEN_2886; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2888 = 12'hb48 == io_in ? 12'hfa1 : _GEN_2887; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2889 = 12'hb49 == io_in ? 12'h24b : _GEN_2888; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2890 = 12'hb4a == io_in ? 12'ha24 : _GEN_2889; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2891 = 12'hb4b == io_in ? 12'h486 : _GEN_2890; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2892 = 12'hb4c == io_in ? 12'h673 : _GEN_2891; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2893 = 12'hb4d == io_in ? 12'h73d : _GEN_2892; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2894 = 12'hb4e == io_in ? 12'h1c7 : _GEN_2893; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2895 = 12'hb4f == io_in ? 12'h26 : _GEN_2894; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2896 = 12'hb50 == io_in ? 12'h26a : _GEN_2895; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2897 = 12'hb51 == io_in ? 12'hddf : _GEN_2896; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2898 = 12'hb52 == io_in ? 12'hcfc : _GEN_2897; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2899 = 12'hb53 == io_in ? 12'h37d : _GEN_2898; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2900 = 12'hb54 == io_in ? 12'hb24 : _GEN_2899; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2901 = 12'hb55 == io_in ? 12'h9d4 : _GEN_2900; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2902 = 12'hb56 == io_in ? 12'he44 : _GEN_2901; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2903 = 12'hb57 == io_in ? 12'hfbf : _GEN_2902; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2904 = 12'hb58 == io_in ? 12'h80f : _GEN_2903; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2905 = 12'hb59 == io_in ? 12'h204 : _GEN_2904; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2906 = 12'hb5a == io_in ? 12'h52a : _GEN_2905; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2907 = 12'hb5b == io_in ? 12'hdad : _GEN_2906; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2908 = 12'hb5c == io_in ? 12'h66f : _GEN_2907; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2909 = 12'hb5d == io_in ? 12'h8a8 : _GEN_2908; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2910 = 12'hb5e == io_in ? 12'h7a2 : _GEN_2909; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2911 = 12'hb5f == io_in ? 12'hf04 : _GEN_2910; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2912 = 12'hb60 == io_in ? 12'hfb1 : _GEN_2911; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2913 = 12'hb61 == io_in ? 12'h478 : _GEN_2912; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2914 = 12'hb62 == io_in ? 12'h206 : _GEN_2913; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2915 = 12'hb63 == io_in ? 12'h9c6 : _GEN_2914; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2916 = 12'hb64 == io_in ? 12'h306 : _GEN_2915; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2917 = 12'hb65 == io_in ? 12'h174 : _GEN_2916; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2918 = 12'hb66 == io_in ? 12'h6dc : _GEN_2917; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2919 = 12'hb67 == io_in ? 12'hb76 : _GEN_2918; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2920 = 12'hb68 == io_in ? 12'h51b : _GEN_2919; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2921 = 12'hb69 == io_in ? 12'h513 : _GEN_2920; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2922 = 12'hb6a == io_in ? 12'he1e : _GEN_2921; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2923 = 12'hb6b == io_in ? 12'h2e1 : _GEN_2922; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2924 = 12'hb6c == io_in ? 12'h914 : _GEN_2923; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2925 = 12'hb6d == io_in ? 12'hd94 : _GEN_2924; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2926 = 12'hb6e == io_in ? 12'h5bb : _GEN_2925; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2927 = 12'hb6f == io_in ? 12'h18d : _GEN_2926; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2928 = 12'hb70 == io_in ? 12'h6eb : _GEN_2927; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2929 = 12'hb71 == io_in ? 12'h1ab : _GEN_2928; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2930 = 12'hb72 == io_in ? 12'h8db : _GEN_2929; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2931 = 12'hb73 == io_in ? 12'h46b : _GEN_2930; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2932 = 12'hb74 == io_in ? 12'h683 : _GEN_2931; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2933 = 12'hb75 == io_in ? 12'he96 : _GEN_2932; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2934 = 12'hb76 == io_in ? 12'ha9 : _GEN_2933; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2935 = 12'hb77 == io_in ? 12'hfb3 : _GEN_2934; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2936 = 12'hb78 == io_in ? 12'hefa : _GEN_2935; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2937 = 12'hb79 == io_in ? 12'h221 : _GEN_2936; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2938 = 12'hb7a == io_in ? 12'h4dd : _GEN_2937; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2939 = 12'hb7b == io_in ? 12'h261 : _GEN_2938; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2940 = 12'hb7c == io_in ? 12'h27a : _GEN_2939; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2941 = 12'hb7d == io_in ? 12'h633 : _GEN_2940; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2942 = 12'hb7e == io_in ? 12'h1cb : _GEN_2941; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2943 = 12'hb7f == io_in ? 12'h907 : _GEN_2942; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2944 = 12'hb80 == io_in ? 12'he13 : _GEN_2943; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2945 = 12'hb81 == io_in ? 12'h87 : _GEN_2944; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2946 = 12'hb82 == io_in ? 12'h93e : _GEN_2945; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2947 = 12'hb83 == io_in ? 12'h841 : _GEN_2946; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2948 = 12'hb84 == io_in ? 12'h41 : _GEN_2947; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2949 = 12'hb85 == io_in ? 12'h520 : _GEN_2948; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2950 = 12'hb86 == io_in ? 12'h6c5 : _GEN_2949; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2951 = 12'hb87 == io_in ? 12'h51 : _GEN_2950; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2952 = 12'hb88 == io_in ? 12'h8dc : _GEN_2951; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2953 = 12'hb89 == io_in ? 12'h23e : _GEN_2952; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2954 = 12'hb8a == io_in ? 12'h1a9 : _GEN_2953; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2955 = 12'hb8b == io_in ? 12'h440 : _GEN_2954; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2956 = 12'hb8c == io_in ? 12'h99d : _GEN_2955; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2957 = 12'hb8d == io_in ? 12'h2e4 : _GEN_2956; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2958 = 12'hb8e == io_in ? 12'h96e : _GEN_2957; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2959 = 12'hb8f == io_in ? 12'hefa : _GEN_2958; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2960 = 12'hb90 == io_in ? 12'h2e4 : _GEN_2959; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2961 = 12'hb91 == io_in ? 12'h7d3 : _GEN_2960; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2962 = 12'hb92 == io_in ? 12'hdb1 : _GEN_2961; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2963 = 12'hb93 == io_in ? 12'h418 : _GEN_2962; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2964 = 12'hb94 == io_in ? 12'h734 : _GEN_2963; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2965 = 12'hb95 == io_in ? 12'h5a : _GEN_2964; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2966 = 12'hb96 == io_in ? 12'h96e : _GEN_2965; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2967 = 12'hb97 == io_in ? 12'h40d : _GEN_2966; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2968 = 12'hb98 == io_in ? 12'h689 : _GEN_2967; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2969 = 12'hb99 == io_in ? 12'hb22 : _GEN_2968; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2970 = 12'hb9a == io_in ? 12'ha77 : _GEN_2969; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2971 = 12'hb9b == io_in ? 12'hd21 : _GEN_2970; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2972 = 12'hb9c == io_in ? 12'h673 : _GEN_2971; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2973 = 12'hb9d == io_in ? 12'he64 : _GEN_2972; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2974 = 12'hb9e == io_in ? 12'h8be : _GEN_2973; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2975 = 12'hb9f == io_in ? 12'hba6 : _GEN_2974; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2976 = 12'hba0 == io_in ? 12'hcbd : _GEN_2975; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2977 = 12'hba1 == io_in ? 12'h56a : _GEN_2976; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2978 = 12'hba2 == io_in ? 12'h332 : _GEN_2977; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2979 = 12'hba3 == io_in ? 12'h201 : _GEN_2978; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2980 = 12'hba4 == io_in ? 12'hff9 : _GEN_2979; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2981 = 12'hba5 == io_in ? 12'h2ae : _GEN_2980; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2982 = 12'hba6 == io_in ? 12'hfa5 : _GEN_2981; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2983 = 12'hba7 == io_in ? 12'h44 : _GEN_2982; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2984 = 12'hba8 == io_in ? 12'he1b : _GEN_2983; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2985 = 12'hba9 == io_in ? 12'h99c : _GEN_2984; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2986 = 12'hbaa == io_in ? 12'hcd6 : _GEN_2985; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2987 = 12'hbab == io_in ? 12'h5b0 : _GEN_2986; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2988 = 12'hbac == io_in ? 12'hf5b : _GEN_2987; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2989 = 12'hbad == io_in ? 12'hd5c : _GEN_2988; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2990 = 12'hbae == io_in ? 12'hddc : _GEN_2989; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2991 = 12'hbaf == io_in ? 12'h4fc : _GEN_2990; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2992 = 12'hbb0 == io_in ? 12'h51 : _GEN_2991; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2993 = 12'hbb1 == io_in ? 12'h24b : _GEN_2992; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2994 = 12'hbb2 == io_in ? 12'hf85 : _GEN_2993; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2995 = 12'hbb3 == io_in ? 12'hd24 : _GEN_2994; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2996 = 12'hbb4 == io_in ? 12'h5b1 : _GEN_2995; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2997 = 12'hbb5 == io_in ? 12'h3c5 : _GEN_2996; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2998 = 12'hbb6 == io_in ? 12'he14 : _GEN_2997; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_2999 = 12'hbb7 == io_in ? 12'h185 : _GEN_2998; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3000 = 12'hbb8 == io_in ? 12'he38 : _GEN_2999; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3001 = 12'hbb9 == io_in ? 12'h656 : _GEN_3000; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3002 = 12'hbba == io_in ? 12'h544 : _GEN_3001; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3003 = 12'hbbb == io_in ? 12'h76d : _GEN_3002; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3004 = 12'hbbc == io_in ? 12'h333 : _GEN_3003; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3005 = 12'hbbd == io_in ? 12'he58 : _GEN_3004; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3006 = 12'hbbe == io_in ? 12'hf31 : _GEN_3005; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3007 = 12'hbbf == io_in ? 12'hfa6 : _GEN_3006; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3008 = 12'hbc0 == io_in ? 12'h779 : _GEN_3007; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3009 = 12'hbc1 == io_in ? 12'hb82 : _GEN_3008; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3010 = 12'hbc2 == io_in ? 12'hbf : _GEN_3009; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3011 = 12'hbc3 == io_in ? 12'hea0 : _GEN_3010; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3012 = 12'hbc4 == io_in ? 12'h1aa : _GEN_3011; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3013 = 12'hbc5 == io_in ? 12'ha1f : _GEN_3012; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3014 = 12'hbc6 == io_in ? 12'h320 : _GEN_3013; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3015 = 12'hbc7 == io_in ? 12'hc7f : _GEN_3014; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3016 = 12'hbc8 == io_in ? 12'h513 : _GEN_3015; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3017 = 12'hbc9 == io_in ? 12'h2dc : _GEN_3016; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3018 = 12'hbca == io_in ? 12'hb3 : _GEN_3017; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3019 = 12'hbcb == io_in ? 12'h352 : _GEN_3018; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3020 = 12'hbcc == io_in ? 12'h172 : _GEN_3019; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3021 = 12'hbcd == io_in ? 12'h93a : _GEN_3020; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3022 = 12'hbce == io_in ? 12'he3f : _GEN_3021; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3023 = 12'hbcf == io_in ? 12'hfbf : _GEN_3022; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3024 = 12'hbd0 == io_in ? 12'h374 : _GEN_3023; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3025 = 12'hbd1 == io_in ? 12'hfe4 : _GEN_3024; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3026 = 12'hbd2 == io_in ? 12'hd01 : _GEN_3025; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3027 = 12'hbd3 == io_in ? 12'h81f : _GEN_3026; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3028 = 12'hbd4 == io_in ? 12'hd34 : _GEN_3027; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3029 = 12'hbd5 == io_in ? 12'h11f : _GEN_3028; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3030 = 12'hbd6 == io_in ? 12'hbec : _GEN_3029; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3031 = 12'hbd7 == io_in ? 12'h6d6 : _GEN_3030; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3032 = 12'hbd8 == io_in ? 12'h87d : _GEN_3031; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3033 = 12'hbd9 == io_in ? 12'h11b : _GEN_3032; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3034 = 12'hbda == io_in ? 12'h921 : _GEN_3033; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3035 = 12'hbdb == io_in ? 12'haf3 : _GEN_3034; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3036 = 12'hbdc == io_in ? 12'h584 : _GEN_3035; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3037 = 12'hbdd == io_in ? 12'h12f : _GEN_3036; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3038 = 12'hbde == io_in ? 12'h4d0 : _GEN_3037; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3039 = 12'hbdf == io_in ? 12'haae : _GEN_3038; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3040 = 12'hbe0 == io_in ? 12'h3e7 : _GEN_3039; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3041 = 12'hbe1 == io_in ? 12'h6c7 : _GEN_3040; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3042 = 12'hbe2 == io_in ? 12'hd1c : _GEN_3041; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3043 = 12'hbe3 == io_in ? 12'h6a1 : _GEN_3042; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3044 = 12'hbe4 == io_in ? 12'hce3 : _GEN_3043; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3045 = 12'hbe5 == io_in ? 12'hb8 : _GEN_3044; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3046 = 12'hbe6 == io_in ? 12'ha29 : _GEN_3045; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3047 = 12'hbe7 == io_in ? 12'hb7e : _GEN_3046; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3048 = 12'hbe8 == io_in ? 12'h367 : _GEN_3047; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3049 = 12'hbe9 == io_in ? 12'hb4a : _GEN_3048; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3050 = 12'hbea == io_in ? 12'h200 : _GEN_3049; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3051 = 12'hbeb == io_in ? 12'h891 : _GEN_3050; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3052 = 12'hbec == io_in ? 12'hec9 : _GEN_3051; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3053 = 12'hbed == io_in ? 12'h4c : _GEN_3052; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3054 = 12'hbee == io_in ? 12'he54 : _GEN_3053; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3055 = 12'hbef == io_in ? 12'hfd9 : _GEN_3054; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3056 = 12'hbf0 == io_in ? 12'he9 : _GEN_3055; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3057 = 12'hbf1 == io_in ? 12'h7a9 : _GEN_3056; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3058 = 12'hbf2 == io_in ? 12'hfa : _GEN_3057; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3059 = 12'hbf3 == io_in ? 12'hc05 : _GEN_3058; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3060 = 12'hbf4 == io_in ? 12'h896 : _GEN_3059; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3061 = 12'hbf5 == io_in ? 12'hfb4 : _GEN_3060; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3062 = 12'hbf6 == io_in ? 12'h674 : _GEN_3061; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3063 = 12'hbf7 == io_in ? 12'h215 : _GEN_3062; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3064 = 12'hbf8 == io_in ? 12'h114 : _GEN_3063; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3065 = 12'hbf9 == io_in ? 12'h660 : _GEN_3064; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3066 = 12'hbfa == io_in ? 12'hd51 : _GEN_3065; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3067 = 12'hbfb == io_in ? 12'h6cd : _GEN_3066; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3068 = 12'hbfc == io_in ? 12'h278 : _GEN_3067; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3069 = 12'hbfd == io_in ? 12'h7c9 : _GEN_3068; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3070 = 12'hbfe == io_in ? 12'h334 : _GEN_3069; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3071 = 12'hbff == io_in ? 12'h19b : _GEN_3070; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3072 = 12'hc00 == io_in ? 12'ha76 : _GEN_3071; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3073 = 12'hc01 == io_in ? 12'hef3 : _GEN_3072; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3074 = 12'hc02 == io_in ? 12'h91 : _GEN_3073; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3075 = 12'hc03 == io_in ? 12'h1fb : _GEN_3074; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3076 = 12'hc04 == io_in ? 12'h792 : _GEN_3075; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3077 = 12'hc05 == io_in ? 12'hdae : _GEN_3076; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3078 = 12'hc06 == io_in ? 12'hf17 : _GEN_3077; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3079 = 12'hc07 == io_in ? 12'h4e4 : _GEN_3078; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3080 = 12'hc08 == io_in ? 12'h256 : _GEN_3079; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3081 = 12'hc09 == io_in ? 12'hd1e : _GEN_3080; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3082 = 12'hc0a == io_in ? 12'h630 : _GEN_3081; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3083 = 12'hc0b == io_in ? 12'hc6d : _GEN_3082; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3084 = 12'hc0c == io_in ? 12'h8c7 : _GEN_3083; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3085 = 12'hc0d == io_in ? 12'h3ff : _GEN_3084; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3086 = 12'hc0e == io_in ? 12'hfff : _GEN_3085; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3087 = 12'hc0f == io_in ? 12'hc29 : _GEN_3086; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3088 = 12'hc10 == io_in ? 12'h388 : _GEN_3087; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3089 = 12'hc11 == io_in ? 12'hfd2 : _GEN_3088; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3090 = 12'hc12 == io_in ? 12'h45 : _GEN_3089; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3091 = 12'hc13 == io_in ? 12'hccd : _GEN_3090; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3092 = 12'hc14 == io_in ? 12'hbff : _GEN_3091; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3093 = 12'hc15 == io_in ? 12'h5ce : _GEN_3092; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3094 = 12'hc16 == io_in ? 12'h70c : _GEN_3093; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3095 = 12'hc17 == io_in ? 12'h50c : _GEN_3094; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3096 = 12'hc18 == io_in ? 12'hd1f : _GEN_3095; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3097 = 12'hc19 == io_in ? 12'h5bd : _GEN_3096; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3098 = 12'hc1a == io_in ? 12'h1ae : _GEN_3097; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3099 = 12'hc1b == io_in ? 12'h4da : _GEN_3098; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3100 = 12'hc1c == io_in ? 12'ha90 : _GEN_3099; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3101 = 12'hc1d == io_in ? 12'h729 : _GEN_3100; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3102 = 12'hc1e == io_in ? 12'h627 : _GEN_3101; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3103 = 12'hc1f == io_in ? 12'hbe6 : _GEN_3102; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3104 = 12'hc20 == io_in ? 12'h338 : _GEN_3103; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3105 = 12'hc21 == io_in ? 12'h73f : _GEN_3104; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3106 = 12'hc22 == io_in ? 12'h36e : _GEN_3105; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3107 = 12'hc23 == io_in ? 12'h8ae : _GEN_3106; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3108 = 12'hc24 == io_in ? 12'hd19 : _GEN_3107; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3109 = 12'hc25 == io_in ? 12'hf5e : _GEN_3108; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3110 = 12'hc26 == io_in ? 12'hcf5 : _GEN_3109; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3111 = 12'hc27 == io_in ? 12'h64 : _GEN_3110; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3112 = 12'hc28 == io_in ? 12'habd : _GEN_3111; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3113 = 12'hc29 == io_in ? 12'h85a : _GEN_3112; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3114 = 12'hc2a == io_in ? 12'hac2 : _GEN_3113; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3115 = 12'hc2b == io_in ? 12'h1da : _GEN_3114; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3116 = 12'hc2c == io_in ? 12'h8e1 : _GEN_3115; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3117 = 12'hc2d == io_in ? 12'h203 : _GEN_3116; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3118 = 12'hc2e == io_in ? 12'h836 : _GEN_3117; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3119 = 12'hc2f == io_in ? 12'h8be : _GEN_3118; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3120 = 12'hc30 == io_in ? 12'ha25 : _GEN_3119; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3121 = 12'hc31 == io_in ? 12'h84a : _GEN_3120; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3122 = 12'hc32 == io_in ? 12'hbe4 : _GEN_3121; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3123 = 12'hc33 == io_in ? 12'h9 : _GEN_3122; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3124 = 12'hc34 == io_in ? 12'h366 : _GEN_3123; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3125 = 12'hc35 == io_in ? 12'h534 : _GEN_3124; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3126 = 12'hc36 == io_in ? 12'h5f7 : _GEN_3125; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3127 = 12'hc37 == io_in ? 12'hb2 : _GEN_3126; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3128 = 12'hc38 == io_in ? 12'hd0b : _GEN_3127; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3129 = 12'hc39 == io_in ? 12'h1a : _GEN_3128; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3130 = 12'hc3a == io_in ? 12'h222 : _GEN_3129; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3131 = 12'hc3b == io_in ? 12'h71c : _GEN_3130; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3132 = 12'hc3c == io_in ? 12'hbaa : _GEN_3131; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3133 = 12'hc3d == io_in ? 12'h555 : _GEN_3132; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3134 = 12'hc3e == io_in ? 12'h73a : _GEN_3133; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3135 = 12'hc3f == io_in ? 12'h16 : _GEN_3134; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3136 = 12'hc40 == io_in ? 12'he82 : _GEN_3135; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3137 = 12'hc41 == io_in ? 12'hdaa : _GEN_3136; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3138 = 12'hc42 == io_in ? 12'h960 : _GEN_3137; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3139 = 12'hc43 == io_in ? 12'hd6a : _GEN_3138; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3140 = 12'hc44 == io_in ? 12'he3b : _GEN_3139; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3141 = 12'hc45 == io_in ? 12'h11c : _GEN_3140; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3142 = 12'hc46 == io_in ? 12'hc31 : _GEN_3141; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3143 = 12'hc47 == io_in ? 12'hfb7 : _GEN_3142; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3144 = 12'hc48 == io_in ? 12'h6e8 : _GEN_3143; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3145 = 12'hc49 == io_in ? 12'h538 : _GEN_3144; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3146 = 12'hc4a == io_in ? 12'hedd : _GEN_3145; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3147 = 12'hc4b == io_in ? 12'h425 : _GEN_3146; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3148 = 12'hc4c == io_in ? 12'h8f3 : _GEN_3147; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3149 = 12'hc4d == io_in ? 12'hb74 : _GEN_3148; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3150 = 12'hc4e == io_in ? 12'hb41 : _GEN_3149; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3151 = 12'hc4f == io_in ? 12'hadb : _GEN_3150; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3152 = 12'hc50 == io_in ? 12'h50e : _GEN_3151; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3153 = 12'hc51 == io_in ? 12'hbb : _GEN_3152; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3154 = 12'hc52 == io_in ? 12'hf78 : _GEN_3153; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3155 = 12'hc53 == io_in ? 12'hf94 : _GEN_3154; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3156 = 12'hc54 == io_in ? 12'hde6 : _GEN_3155; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3157 = 12'hc55 == io_in ? 12'hc3d : _GEN_3156; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3158 = 12'hc56 == io_in ? 12'h4ab : _GEN_3157; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3159 = 12'hc57 == io_in ? 12'hfa9 : _GEN_3158; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3160 = 12'hc58 == io_in ? 12'h84c : _GEN_3159; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3161 = 12'hc59 == io_in ? 12'h1e4 : _GEN_3160; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3162 = 12'hc5a == io_in ? 12'h72 : _GEN_3161; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3163 = 12'hc5b == io_in ? 12'h52c : _GEN_3162; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3164 = 12'hc5c == io_in ? 12'h9cd : _GEN_3163; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3165 = 12'hc5d == io_in ? 12'hcd1 : _GEN_3164; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3166 = 12'hc5e == io_in ? 12'h4ad : _GEN_3165; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3167 = 12'hc5f == io_in ? 12'h14c : _GEN_3166; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3168 = 12'hc60 == io_in ? 12'h153 : _GEN_3167; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3169 = 12'hc61 == io_in ? 12'h9d5 : _GEN_3168; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3170 = 12'hc62 == io_in ? 12'hd10 : _GEN_3169; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3171 = 12'hc63 == io_in ? 12'ha46 : _GEN_3170; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3172 = 12'hc64 == io_in ? 12'h1cf : _GEN_3171; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3173 = 12'hc65 == io_in ? 12'h98f : _GEN_3172; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3174 = 12'hc66 == io_in ? 12'h491 : _GEN_3173; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3175 = 12'hc67 == io_in ? 12'hbaa : _GEN_3174; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3176 = 12'hc68 == io_in ? 12'h238 : _GEN_3175; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3177 = 12'hc69 == io_in ? 12'h829 : _GEN_3176; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3178 = 12'hc6a == io_in ? 12'h74b : _GEN_3177; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3179 = 12'hc6b == io_in ? 12'h776 : _GEN_3178; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3180 = 12'hc6c == io_in ? 12'h670 : _GEN_3179; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3181 = 12'hc6d == io_in ? 12'h69f : _GEN_3180; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3182 = 12'hc6e == io_in ? 12'h842 : _GEN_3181; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3183 = 12'hc6f == io_in ? 12'h201 : _GEN_3182; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3184 = 12'hc70 == io_in ? 12'hb67 : _GEN_3183; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3185 = 12'hc71 == io_in ? 12'h235 : _GEN_3184; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3186 = 12'hc72 == io_in ? 12'h40d : _GEN_3185; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3187 = 12'hc73 == io_in ? 12'h253 : _GEN_3186; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3188 = 12'hc74 == io_in ? 12'hdd8 : _GEN_3187; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3189 = 12'hc75 == io_in ? 12'h37a : _GEN_3188; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3190 = 12'hc76 == io_in ? 12'h175 : _GEN_3189; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3191 = 12'hc77 == io_in ? 12'h7cc : _GEN_3190; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3192 = 12'hc78 == io_in ? 12'hae9 : _GEN_3191; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3193 = 12'hc79 == io_in ? 12'h2d2 : _GEN_3192; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3194 = 12'hc7a == io_in ? 12'hc5b : _GEN_3193; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3195 = 12'hc7b == io_in ? 12'h1c2 : _GEN_3194; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3196 = 12'hc7c == io_in ? 12'h6b7 : _GEN_3195; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3197 = 12'hc7d == io_in ? 12'hea8 : _GEN_3196; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3198 = 12'hc7e == io_in ? 12'hba1 : _GEN_3197; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3199 = 12'hc7f == io_in ? 12'h5cf : _GEN_3198; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3200 = 12'hc80 == io_in ? 12'hd9a : _GEN_3199; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3201 = 12'hc81 == io_in ? 12'h36a : _GEN_3200; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3202 = 12'hc82 == io_in ? 12'h412 : _GEN_3201; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3203 = 12'hc83 == io_in ? 12'h789 : _GEN_3202; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3204 = 12'hc84 == io_in ? 12'he50 : _GEN_3203; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3205 = 12'hc85 == io_in ? 12'h99d : _GEN_3204; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3206 = 12'hc86 == io_in ? 12'hc84 : _GEN_3205; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3207 = 12'hc87 == io_in ? 12'hc31 : _GEN_3206; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3208 = 12'hc88 == io_in ? 12'he90 : _GEN_3207; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3209 = 12'hc89 == io_in ? 12'hf63 : _GEN_3208; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3210 = 12'hc8a == io_in ? 12'h4b7 : _GEN_3209; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3211 = 12'hc8b == io_in ? 12'h556 : _GEN_3210; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3212 = 12'hc8c == io_in ? 12'h85e : _GEN_3211; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3213 = 12'hc8d == io_in ? 12'h355 : _GEN_3212; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3214 = 12'hc8e == io_in ? 12'hc1a : _GEN_3213; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3215 = 12'hc8f == io_in ? 12'he0a : _GEN_3214; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3216 = 12'hc90 == io_in ? 12'h4c : _GEN_3215; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3217 = 12'hc91 == io_in ? 12'h45f : _GEN_3216; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3218 = 12'hc92 == io_in ? 12'hf2d : _GEN_3217; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3219 = 12'hc93 == io_in ? 12'h304 : _GEN_3218; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3220 = 12'hc94 == io_in ? 12'h5cb : _GEN_3219; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3221 = 12'hc95 == io_in ? 12'hfe5 : _GEN_3220; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3222 = 12'hc96 == io_in ? 12'hc67 : _GEN_3221; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3223 = 12'hc97 == io_in ? 12'had5 : _GEN_3222; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3224 = 12'hc98 == io_in ? 12'hcd7 : _GEN_3223; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3225 = 12'hc99 == io_in ? 12'h33e : _GEN_3224; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3226 = 12'hc9a == io_in ? 12'h1fc : _GEN_3225; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3227 = 12'hc9b == io_in ? 12'h40 : _GEN_3226; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3228 = 12'hc9c == io_in ? 12'h47 : _GEN_3227; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3229 = 12'hc9d == io_in ? 12'hb05 : _GEN_3228; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3230 = 12'hc9e == io_in ? 12'hd9e : _GEN_3229; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3231 = 12'hc9f == io_in ? 12'heba : _GEN_3230; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3232 = 12'hca0 == io_in ? 12'he42 : _GEN_3231; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3233 = 12'hca1 == io_in ? 12'h81b : _GEN_3232; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3234 = 12'hca2 == io_in ? 12'h324 : _GEN_3233; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3235 = 12'hca3 == io_in ? 12'h47d : _GEN_3234; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3236 = 12'hca4 == io_in ? 12'h42e : _GEN_3235; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3237 = 12'hca5 == io_in ? 12'h3e7 : _GEN_3236; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3238 = 12'hca6 == io_in ? 12'hdb3 : _GEN_3237; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3239 = 12'hca7 == io_in ? 12'h397 : _GEN_3238; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3240 = 12'hca8 == io_in ? 12'h79e : _GEN_3239; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3241 = 12'hca9 == io_in ? 12'h1fc : _GEN_3240; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3242 = 12'hcaa == io_in ? 12'h445 : _GEN_3241; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3243 = 12'hcab == io_in ? 12'hd4d : _GEN_3242; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3244 = 12'hcac == io_in ? 12'h21 : _GEN_3243; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3245 = 12'hcad == io_in ? 12'h9c1 : _GEN_3244; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3246 = 12'hcae == io_in ? 12'h391 : _GEN_3245; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3247 = 12'hcaf == io_in ? 12'ha5b : _GEN_3246; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3248 = 12'hcb0 == io_in ? 12'hfcd : _GEN_3247; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3249 = 12'hcb1 == io_in ? 12'h637 : _GEN_3248; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3250 = 12'hcb2 == io_in ? 12'h64e : _GEN_3249; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3251 = 12'hcb3 == io_in ? 12'hd1a : _GEN_3250; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3252 = 12'hcb4 == io_in ? 12'ha3d : _GEN_3251; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3253 = 12'hcb5 == io_in ? 12'h1a8 : _GEN_3252; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3254 = 12'hcb6 == io_in ? 12'h59f : _GEN_3253; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3255 = 12'hcb7 == io_in ? 12'he0d : _GEN_3254; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3256 = 12'hcb8 == io_in ? 12'hb21 : _GEN_3255; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3257 = 12'hcb9 == io_in ? 12'hf09 : _GEN_3256; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3258 = 12'hcba == io_in ? 12'h695 : _GEN_3257; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3259 = 12'hcbb == io_in ? 12'h25d : _GEN_3258; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3260 = 12'hcbc == io_in ? 12'hdaf : _GEN_3259; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3261 = 12'hcbd == io_in ? 12'h856 : _GEN_3260; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3262 = 12'hcbe == io_in ? 12'h96c : _GEN_3261; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3263 = 12'hcbf == io_in ? 12'h8aa : _GEN_3262; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3264 = 12'hcc0 == io_in ? 12'hf10 : _GEN_3263; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3265 = 12'hcc1 == io_in ? 12'h928 : _GEN_3264; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3266 = 12'hcc2 == io_in ? 12'habd : _GEN_3265; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3267 = 12'hcc3 == io_in ? 12'ha5b : _GEN_3266; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3268 = 12'hcc4 == io_in ? 12'hfb : _GEN_3267; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3269 = 12'hcc5 == io_in ? 12'h4d3 : _GEN_3268; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3270 = 12'hcc6 == io_in ? 12'h6f1 : _GEN_3269; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3271 = 12'hcc7 == io_in ? 12'h4b4 : _GEN_3270; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3272 = 12'hcc8 == io_in ? 12'hbeb : _GEN_3271; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3273 = 12'hcc9 == io_in ? 12'h89c : _GEN_3272; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3274 = 12'hcca == io_in ? 12'h272 : _GEN_3273; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3275 = 12'hccb == io_in ? 12'h18b : _GEN_3274; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3276 = 12'hccc == io_in ? 12'hd19 : _GEN_3275; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3277 = 12'hccd == io_in ? 12'hbe5 : _GEN_3276; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3278 = 12'hcce == io_in ? 12'h4d7 : _GEN_3277; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3279 = 12'hccf == io_in ? 12'h61d : _GEN_3278; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3280 = 12'hcd0 == io_in ? 12'hbb1 : _GEN_3279; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3281 = 12'hcd1 == io_in ? 12'h266 : _GEN_3280; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3282 = 12'hcd2 == io_in ? 12'he83 : _GEN_3281; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3283 = 12'hcd3 == io_in ? 12'h7ae : _GEN_3282; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3284 = 12'hcd4 == io_in ? 12'h31 : _GEN_3283; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3285 = 12'hcd5 == io_in ? 12'h770 : _GEN_3284; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3286 = 12'hcd6 == io_in ? 12'hcd3 : _GEN_3285; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3287 = 12'hcd7 == io_in ? 12'h10b : _GEN_3286; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3288 = 12'hcd8 == io_in ? 12'hae3 : _GEN_3287; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3289 = 12'hcd9 == io_in ? 12'he12 : _GEN_3288; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3290 = 12'hcda == io_in ? 12'hb8f : _GEN_3289; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3291 = 12'hcdb == io_in ? 12'h5d2 : _GEN_3290; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3292 = 12'hcdc == io_in ? 12'h379 : _GEN_3291; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3293 = 12'hcdd == io_in ? 12'h109 : _GEN_3292; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3294 = 12'hcde == io_in ? 12'hf36 : _GEN_3293; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3295 = 12'hcdf == io_in ? 12'hd88 : _GEN_3294; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3296 = 12'hce0 == io_in ? 12'h852 : _GEN_3295; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3297 = 12'hce1 == io_in ? 12'h87d : _GEN_3296; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3298 = 12'hce2 == io_in ? 12'h3f0 : _GEN_3297; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3299 = 12'hce3 == io_in ? 12'h13e : _GEN_3298; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3300 = 12'hce4 == io_in ? 12'h363 : _GEN_3299; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3301 = 12'hce5 == io_in ? 12'h32d : _GEN_3300; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3302 = 12'hce6 == io_in ? 12'h372 : _GEN_3301; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3303 = 12'hce7 == io_in ? 12'hc32 : _GEN_3302; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3304 = 12'hce8 == io_in ? 12'h3bb : _GEN_3303; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3305 = 12'hce9 == io_in ? 12'h7bb : _GEN_3304; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3306 = 12'hcea == io_in ? 12'h84a : _GEN_3305; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3307 = 12'hceb == io_in ? 12'h7a4 : _GEN_3306; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3308 = 12'hcec == io_in ? 12'hb0f : _GEN_3307; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3309 = 12'hced == io_in ? 12'h18f : _GEN_3308; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3310 = 12'hcee == io_in ? 12'h850 : _GEN_3309; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3311 = 12'hcef == io_in ? 12'h18d : _GEN_3310; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3312 = 12'hcf0 == io_in ? 12'he : _GEN_3311; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3313 = 12'hcf1 == io_in ? 12'h723 : _GEN_3312; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3314 = 12'hcf2 == io_in ? 12'h89 : _GEN_3313; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3315 = 12'hcf3 == io_in ? 12'h683 : _GEN_3314; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3316 = 12'hcf4 == io_in ? 12'h8e : _GEN_3315; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3317 = 12'hcf5 == io_in ? 12'he50 : _GEN_3316; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3318 = 12'hcf6 == io_in ? 12'ha36 : _GEN_3317; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3319 = 12'hcf7 == io_in ? 12'hb87 : _GEN_3318; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3320 = 12'hcf8 == io_in ? 12'he18 : _GEN_3319; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3321 = 12'hcf9 == io_in ? 12'ha3a : _GEN_3320; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3322 = 12'hcfa == io_in ? 12'hfd9 : _GEN_3321; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3323 = 12'hcfb == io_in ? 12'ha21 : _GEN_3322; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3324 = 12'hcfc == io_in ? 12'h65b : _GEN_3323; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3325 = 12'hcfd == io_in ? 12'hfd5 : _GEN_3324; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3326 = 12'hcfe == io_in ? 12'h800 : _GEN_3325; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3327 = 12'hcff == io_in ? 12'hf5b : _GEN_3326; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3328 = 12'hd00 == io_in ? 12'h65f : _GEN_3327; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3329 = 12'hd01 == io_in ? 12'hd57 : _GEN_3328; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3330 = 12'hd02 == io_in ? 12'h598 : _GEN_3329; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3331 = 12'hd03 == io_in ? 12'hf2f : _GEN_3330; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3332 = 12'hd04 == io_in ? 12'h7f5 : _GEN_3331; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3333 = 12'hd05 == io_in ? 12'h14f : _GEN_3332; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3334 = 12'hd06 == io_in ? 12'hf55 : _GEN_3333; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3335 = 12'hd07 == io_in ? 12'h4ee : _GEN_3334; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3336 = 12'hd08 == io_in ? 12'hdc4 : _GEN_3335; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3337 = 12'hd09 == io_in ? 12'h36d : _GEN_3336; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3338 = 12'hd0a == io_in ? 12'haea : _GEN_3337; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3339 = 12'hd0b == io_in ? 12'h55d : _GEN_3338; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3340 = 12'hd0c == io_in ? 12'h371 : _GEN_3339; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3341 = 12'hd0d == io_in ? 12'h6f0 : _GEN_3340; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3342 = 12'hd0e == io_in ? 12'h8af : _GEN_3341; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3343 = 12'hd0f == io_in ? 12'h856 : _GEN_3342; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3344 = 12'hd10 == io_in ? 12'h7ae : _GEN_3343; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3345 = 12'hd11 == io_in ? 12'h9a3 : _GEN_3344; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3346 = 12'hd12 == io_in ? 12'h919 : _GEN_3345; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3347 = 12'hd13 == io_in ? 12'h90a : _GEN_3346; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3348 = 12'hd14 == io_in ? 12'h850 : _GEN_3347; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3349 = 12'hd15 == io_in ? 12'h637 : _GEN_3348; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3350 = 12'hd16 == io_in ? 12'h8a9 : _GEN_3349; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3351 = 12'hd17 == io_in ? 12'ha3a : _GEN_3350; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3352 = 12'hd18 == io_in ? 12'h232 : _GEN_3351; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3353 = 12'hd19 == io_in ? 12'h300 : _GEN_3352; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3354 = 12'hd1a == io_in ? 12'h794 : _GEN_3353; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3355 = 12'hd1b == io_in ? 12'h667 : _GEN_3354; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3356 = 12'hd1c == io_in ? 12'h4dc : _GEN_3355; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3357 = 12'hd1d == io_in ? 12'h28d : _GEN_3356; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3358 = 12'hd1e == io_in ? 12'h86c : _GEN_3357; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3359 = 12'hd1f == io_in ? 12'h42f : _GEN_3358; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3360 = 12'hd20 == io_in ? 12'h4e3 : _GEN_3359; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3361 = 12'hd21 == io_in ? 12'h884 : _GEN_3360; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3362 = 12'hd22 == io_in ? 12'h9d9 : _GEN_3361; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3363 = 12'hd23 == io_in ? 12'h937 : _GEN_3362; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3364 = 12'hd24 == io_in ? 12'h6b9 : _GEN_3363; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3365 = 12'hd25 == io_in ? 12'h6dd : _GEN_3364; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3366 = 12'hd26 == io_in ? 12'h17e : _GEN_3365; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3367 = 12'hd27 == io_in ? 12'hf5b : _GEN_3366; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3368 = 12'hd28 == io_in ? 12'h9ae : _GEN_3367; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3369 = 12'hd29 == io_in ? 12'h4bf : _GEN_3368; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3370 = 12'hd2a == io_in ? 12'h556 : _GEN_3369; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3371 = 12'hd2b == io_in ? 12'h184 : _GEN_3370; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3372 = 12'hd2c == io_in ? 12'h95d : _GEN_3371; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3373 = 12'hd2d == io_in ? 12'h5b9 : _GEN_3372; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3374 = 12'hd2e == io_in ? 12'h26c : _GEN_3373; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3375 = 12'hd2f == io_in ? 12'h103 : _GEN_3374; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3376 = 12'hd30 == io_in ? 12'h847 : _GEN_3375; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3377 = 12'hd31 == io_in ? 12'hd1b : _GEN_3376; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3378 = 12'hd32 == io_in ? 12'hd97 : _GEN_3377; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3379 = 12'hd33 == io_in ? 12'hf8d : _GEN_3378; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3380 = 12'hd34 == io_in ? 12'hd88 : _GEN_3379; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3381 = 12'hd35 == io_in ? 12'h2f4 : _GEN_3380; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3382 = 12'hd36 == io_in ? 12'h93d : _GEN_3381; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3383 = 12'hd37 == io_in ? 12'h2d1 : _GEN_3382; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3384 = 12'hd38 == io_in ? 12'h83 : _GEN_3383; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3385 = 12'hd39 == io_in ? 12'h69f : _GEN_3384; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3386 = 12'hd3a == io_in ? 12'h20e : _GEN_3385; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3387 = 12'hd3b == io_in ? 12'h740 : _GEN_3386; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3388 = 12'hd3c == io_in ? 12'hfcb : _GEN_3387; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3389 = 12'hd3d == io_in ? 12'hb8b : _GEN_3388; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3390 = 12'hd3e == io_in ? 12'h6d1 : _GEN_3389; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3391 = 12'hd3f == io_in ? 12'hb0a : _GEN_3390; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3392 = 12'hd40 == io_in ? 12'h601 : _GEN_3391; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3393 = 12'hd41 == io_in ? 12'h26 : _GEN_3392; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3394 = 12'hd42 == io_in ? 12'hbf2 : _GEN_3393; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3395 = 12'hd43 == io_in ? 12'he87 : _GEN_3394; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3396 = 12'hd44 == io_in ? 12'h99c : _GEN_3395; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3397 = 12'hd45 == io_in ? 12'hb14 : _GEN_3396; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3398 = 12'hd46 == io_in ? 12'h2bd : _GEN_3397; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3399 = 12'hd47 == io_in ? 12'h3ff : _GEN_3398; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3400 = 12'hd48 == io_in ? 12'h866 : _GEN_3399; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3401 = 12'hd49 == io_in ? 12'h8aa : _GEN_3400; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3402 = 12'hd4a == io_in ? 12'h499 : _GEN_3401; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3403 = 12'hd4b == io_in ? 12'hdd : _GEN_3402; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3404 = 12'hd4c == io_in ? 12'h880 : _GEN_3403; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3405 = 12'hd4d == io_in ? 12'hcd : _GEN_3404; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3406 = 12'hd4e == io_in ? 12'ha77 : _GEN_3405; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3407 = 12'hd4f == io_in ? 12'h975 : _GEN_3406; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3408 = 12'hd50 == io_in ? 12'he83 : _GEN_3407; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3409 = 12'hd51 == io_in ? 12'h555 : _GEN_3408; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3410 = 12'hd52 == io_in ? 12'hd01 : _GEN_3409; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3411 = 12'hd53 == io_in ? 12'he57 : _GEN_3410; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3412 = 12'hd54 == io_in ? 12'h12d : _GEN_3411; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3413 = 12'hd55 == io_in ? 12'h1c8 : _GEN_3412; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3414 = 12'hd56 == io_in ? 12'h803 : _GEN_3413; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3415 = 12'hd57 == io_in ? 12'h6eb : _GEN_3414; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3416 = 12'hd58 == io_in ? 12'h87c : _GEN_3415; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3417 = 12'hd59 == io_in ? 12'h8ca : _GEN_3416; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3418 = 12'hd5a == io_in ? 12'h60d : _GEN_3417; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3419 = 12'hd5b == io_in ? 12'hcb6 : _GEN_3418; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3420 = 12'hd5c == io_in ? 12'h97f : _GEN_3419; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3421 = 12'hd5d == io_in ? 12'h9aa : _GEN_3420; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3422 = 12'hd5e == io_in ? 12'hca0 : _GEN_3421; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3423 = 12'hd5f == io_in ? 12'h1f0 : _GEN_3422; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3424 = 12'hd60 == io_in ? 12'hd3d : _GEN_3423; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3425 = 12'hd61 == io_in ? 12'hb15 : _GEN_3424; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3426 = 12'hd62 == io_in ? 12'h656 : _GEN_3425; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3427 = 12'hd63 == io_in ? 12'h5b4 : _GEN_3426; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3428 = 12'hd64 == io_in ? 12'h3a7 : _GEN_3427; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3429 = 12'hd65 == io_in ? 12'h7a6 : _GEN_3428; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3430 = 12'hd66 == io_in ? 12'ha4d : _GEN_3429; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3431 = 12'hd67 == io_in ? 12'h8f8 : _GEN_3430; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3432 = 12'hd68 == io_in ? 12'ha42 : _GEN_3431; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3433 = 12'hd69 == io_in ? 12'h8d : _GEN_3432; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3434 = 12'hd6a == io_in ? 12'he3d : _GEN_3433; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3435 = 12'hd6b == io_in ? 12'h71c : _GEN_3434; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3436 = 12'hd6c == io_in ? 12'hec3 : _GEN_3435; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3437 = 12'hd6d == io_in ? 12'ha7f : _GEN_3436; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3438 = 12'hd6e == io_in ? 12'h44e : _GEN_3437; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3439 = 12'hd6f == io_in ? 12'h877 : _GEN_3438; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3440 = 12'hd70 == io_in ? 12'h1d4 : _GEN_3439; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3441 = 12'hd71 == io_in ? 12'hcd0 : _GEN_3440; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3442 = 12'hd72 == io_in ? 12'h540 : _GEN_3441; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3443 = 12'hd73 == io_in ? 12'h6f4 : _GEN_3442; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3444 = 12'hd74 == io_in ? 12'h5bb : _GEN_3443; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3445 = 12'hd75 == io_in ? 12'hb8e : _GEN_3444; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3446 = 12'hd76 == io_in ? 12'ha30 : _GEN_3445; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3447 = 12'hd77 == io_in ? 12'he2d : _GEN_3446; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3448 = 12'hd78 == io_in ? 12'hbb3 : _GEN_3447; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3449 = 12'hd79 == io_in ? 12'hef0 : _GEN_3448; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3450 = 12'hd7a == io_in ? 12'hc6f : _GEN_3449; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3451 = 12'hd7b == io_in ? 12'h49 : _GEN_3450; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3452 = 12'hd7c == io_in ? 12'h3f0 : _GEN_3451; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3453 = 12'hd7d == io_in ? 12'hecb : _GEN_3452; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3454 = 12'hd7e == io_in ? 12'hb1a : _GEN_3453; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3455 = 12'hd7f == io_in ? 12'h4f8 : _GEN_3454; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3456 = 12'hd80 == io_in ? 12'h640 : _GEN_3455; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3457 = 12'hd81 == io_in ? 12'h3c4 : _GEN_3456; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3458 = 12'hd82 == io_in ? 12'h924 : _GEN_3457; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3459 = 12'hd83 == io_in ? 12'h3f7 : _GEN_3458; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3460 = 12'hd84 == io_in ? 12'h107 : _GEN_3459; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3461 = 12'hd85 == io_in ? 12'hc21 : _GEN_3460; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3462 = 12'hd86 == io_in ? 12'h799 : _GEN_3461; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3463 = 12'hd87 == io_in ? 12'h29a : _GEN_3462; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3464 = 12'hd88 == io_in ? 12'h2f0 : _GEN_3463; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3465 = 12'hd89 == io_in ? 12'hc3c : _GEN_3464; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3466 = 12'hd8a == io_in ? 12'h90a : _GEN_3465; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3467 = 12'hd8b == io_in ? 12'h3f2 : _GEN_3466; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3468 = 12'hd8c == io_in ? 12'h8c6 : _GEN_3467; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3469 = 12'hd8d == io_in ? 12'hd64 : _GEN_3468; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3470 = 12'hd8e == io_in ? 12'hf56 : _GEN_3469; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3471 = 12'hd8f == io_in ? 12'hc59 : _GEN_3470; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3472 = 12'hd90 == io_in ? 12'h81a : _GEN_3471; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3473 = 12'hd91 == io_in ? 12'h672 : _GEN_3472; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3474 = 12'hd92 == io_in ? 12'h4b6 : _GEN_3473; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3475 = 12'hd93 == io_in ? 12'hf82 : _GEN_3474; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3476 = 12'hd94 == io_in ? 12'h2a6 : _GEN_3475; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3477 = 12'hd95 == io_in ? 12'hb6c : _GEN_3476; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3478 = 12'hd96 == io_in ? 12'hd8b : _GEN_3477; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3479 = 12'hd97 == io_in ? 12'hf64 : _GEN_3478; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3480 = 12'hd98 == io_in ? 12'h3c2 : _GEN_3479; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3481 = 12'hd99 == io_in ? 12'ha12 : _GEN_3480; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3482 = 12'hd9a == io_in ? 12'h10d : _GEN_3481; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3483 = 12'hd9b == io_in ? 12'hb02 : _GEN_3482; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3484 = 12'hd9c == io_in ? 12'h599 : _GEN_3483; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3485 = 12'hd9d == io_in ? 12'hcee : _GEN_3484; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3486 = 12'hd9e == io_in ? 12'hb53 : _GEN_3485; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3487 = 12'hd9f == io_in ? 12'he74 : _GEN_3486; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3488 = 12'hda0 == io_in ? 12'hf62 : _GEN_3487; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3489 = 12'hda1 == io_in ? 12'habd : _GEN_3488; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3490 = 12'hda2 == io_in ? 12'he1 : _GEN_3489; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3491 = 12'hda3 == io_in ? 12'h68a : _GEN_3490; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3492 = 12'hda4 == io_in ? 12'h7e9 : _GEN_3491; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3493 = 12'hda5 == io_in ? 12'h9f2 : _GEN_3492; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3494 = 12'hda6 == io_in ? 12'h158 : _GEN_3493; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3495 = 12'hda7 == io_in ? 12'h714 : _GEN_3494; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3496 = 12'hda8 == io_in ? 12'hb3f : _GEN_3495; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3497 = 12'hda9 == io_in ? 12'h5a1 : _GEN_3496; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3498 = 12'hdaa == io_in ? 12'h1e : _GEN_3497; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3499 = 12'hdab == io_in ? 12'h425 : _GEN_3498; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3500 = 12'hdac == io_in ? 12'h92c : _GEN_3499; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3501 = 12'hdad == io_in ? 12'hfb2 : _GEN_3500; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3502 = 12'hdae == io_in ? 12'h38b : _GEN_3501; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3503 = 12'hdaf == io_in ? 12'he99 : _GEN_3502; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3504 = 12'hdb0 == io_in ? 12'h11e : _GEN_3503; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3505 = 12'hdb1 == io_in ? 12'h2c9 : _GEN_3504; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3506 = 12'hdb2 == io_in ? 12'h2e : _GEN_3505; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3507 = 12'hdb3 == io_in ? 12'hf : _GEN_3506; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3508 = 12'hdb4 == io_in ? 12'hc9c : _GEN_3507; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3509 = 12'hdb5 == io_in ? 12'h215 : _GEN_3508; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3510 = 12'hdb6 == io_in ? 12'h134 : _GEN_3509; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3511 = 12'hdb7 == io_in ? 12'hb0 : _GEN_3510; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3512 = 12'hdb8 == io_in ? 12'h9ee : _GEN_3511; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3513 = 12'hdb9 == io_in ? 12'h62b : _GEN_3512; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3514 = 12'hdba == io_in ? 12'h201 : _GEN_3513; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3515 = 12'hdbb == io_in ? 12'h392 : _GEN_3514; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3516 = 12'hdbc == io_in ? 12'hd2d : _GEN_3515; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3517 = 12'hdbd == io_in ? 12'h1db : _GEN_3516; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3518 = 12'hdbe == io_in ? 12'h18e : _GEN_3517; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3519 = 12'hdbf == io_in ? 12'h21 : _GEN_3518; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3520 = 12'hdc0 == io_in ? 12'hd : _GEN_3519; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3521 = 12'hdc1 == io_in ? 12'ha8 : _GEN_3520; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3522 = 12'hdc2 == io_in ? 12'h588 : _GEN_3521; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3523 = 12'hdc3 == io_in ? 12'h60b : _GEN_3522; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3524 = 12'hdc4 == io_in ? 12'h21c : _GEN_3523; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3525 = 12'hdc5 == io_in ? 12'hed : _GEN_3524; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3526 = 12'hdc6 == io_in ? 12'h1f3 : _GEN_3525; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3527 = 12'hdc7 == io_in ? 12'hd2c : _GEN_3526; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3528 = 12'hdc8 == io_in ? 12'h8aa : _GEN_3527; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3529 = 12'hdc9 == io_in ? 12'h5e3 : _GEN_3528; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3530 = 12'hdca == io_in ? 12'h84d : _GEN_3529; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3531 = 12'hdcb == io_in ? 12'hec0 : _GEN_3530; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3532 = 12'hdcc == io_in ? 12'h2b9 : _GEN_3531; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3533 = 12'hdcd == io_in ? 12'h931 : _GEN_3532; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3534 = 12'hdce == io_in ? 12'h57c : _GEN_3533; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3535 = 12'hdcf == io_in ? 12'h4a6 : _GEN_3534; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3536 = 12'hdd0 == io_in ? 12'h1d5 : _GEN_3535; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3537 = 12'hdd1 == io_in ? 12'he2 : _GEN_3536; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3538 = 12'hdd2 == io_in ? 12'h50e : _GEN_3537; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3539 = 12'hdd3 == io_in ? 12'he09 : _GEN_3538; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3540 = 12'hdd4 == io_in ? 12'ha90 : _GEN_3539; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3541 = 12'hdd5 == io_in ? 12'hda5 : _GEN_3540; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3542 = 12'hdd6 == io_in ? 12'hfb0 : _GEN_3541; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3543 = 12'hdd7 == io_in ? 12'h6cd : _GEN_3542; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3544 = 12'hdd8 == io_in ? 12'h8a3 : _GEN_3543; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3545 = 12'hdd9 == io_in ? 12'h724 : _GEN_3544; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3546 = 12'hdda == io_in ? 12'h528 : _GEN_3545; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3547 = 12'hddb == io_in ? 12'hc89 : _GEN_3546; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3548 = 12'hddc == io_in ? 12'hc1d : _GEN_3547; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3549 = 12'hddd == io_in ? 12'h95a : _GEN_3548; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3550 = 12'hdde == io_in ? 12'hbda : _GEN_3549; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3551 = 12'hddf == io_in ? 12'hd71 : _GEN_3550; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3552 = 12'hde0 == io_in ? 12'h2e7 : _GEN_3551; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3553 = 12'hde1 == io_in ? 12'hfec : _GEN_3552; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3554 = 12'hde2 == io_in ? 12'h9ec : _GEN_3553; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3555 = 12'hde3 == io_in ? 12'hbf7 : _GEN_3554; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3556 = 12'hde4 == io_in ? 12'h792 : _GEN_3555; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3557 = 12'hde5 == io_in ? 12'h46a : _GEN_3556; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3558 = 12'hde6 == io_in ? 12'h945 : _GEN_3557; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3559 = 12'hde7 == io_in ? 12'he06 : _GEN_3558; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3560 = 12'hde8 == io_in ? 12'h2c0 : _GEN_3559; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3561 = 12'hde9 == io_in ? 12'hc2d : _GEN_3560; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3562 = 12'hdea == io_in ? 12'hfd8 : _GEN_3561; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3563 = 12'hdeb == io_in ? 12'h649 : _GEN_3562; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3564 = 12'hdec == io_in ? 12'hd3f : _GEN_3563; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3565 = 12'hded == io_in ? 12'h3ba : _GEN_3564; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3566 = 12'hdee == io_in ? 12'h999 : _GEN_3565; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3567 = 12'hdef == io_in ? 12'h5ab : _GEN_3566; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3568 = 12'hdf0 == io_in ? 12'h777 : _GEN_3567; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3569 = 12'hdf1 == io_in ? 12'h2a5 : _GEN_3568; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3570 = 12'hdf2 == io_in ? 12'hfe2 : _GEN_3569; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3571 = 12'hdf3 == io_in ? 12'hdbc : _GEN_3570; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3572 = 12'hdf4 == io_in ? 12'hfa0 : _GEN_3571; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3573 = 12'hdf5 == io_in ? 12'hdfc : _GEN_3572; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3574 = 12'hdf6 == io_in ? 12'h24e : _GEN_3573; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3575 = 12'hdf7 == io_in ? 12'hb5f : _GEN_3574; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3576 = 12'hdf8 == io_in ? 12'hec0 : _GEN_3575; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3577 = 12'hdf9 == io_in ? 12'hb5a : _GEN_3576; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3578 = 12'hdfa == io_in ? 12'hc04 : _GEN_3577; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3579 = 12'hdfb == io_in ? 12'ha96 : _GEN_3578; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3580 = 12'hdfc == io_in ? 12'hfeb : _GEN_3579; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3581 = 12'hdfd == io_in ? 12'hdfa : _GEN_3580; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3582 = 12'hdfe == io_in ? 12'h410 : _GEN_3581; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3583 = 12'hdff == io_in ? 12'hee0 : _GEN_3582; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3584 = 12'he00 == io_in ? 12'hbd3 : _GEN_3583; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3585 = 12'he01 == io_in ? 12'hdd2 : _GEN_3584; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3586 = 12'he02 == io_in ? 12'h367 : _GEN_3585; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3587 = 12'he03 == io_in ? 12'h22d : _GEN_3586; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3588 = 12'he04 == io_in ? 12'h1a0 : _GEN_3587; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3589 = 12'he05 == io_in ? 12'hf1 : _GEN_3588; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3590 = 12'he06 == io_in ? 12'hb9e : _GEN_3589; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3591 = 12'he07 == io_in ? 12'h1fd : _GEN_3590; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3592 = 12'he08 == io_in ? 12'he56 : _GEN_3591; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3593 = 12'he09 == io_in ? 12'hdf6 : _GEN_3592; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3594 = 12'he0a == io_in ? 12'h6c : _GEN_3593; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3595 = 12'he0b == io_in ? 12'h60e : _GEN_3594; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3596 = 12'he0c == io_in ? 12'hd5b : _GEN_3595; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3597 = 12'he0d == io_in ? 12'he49 : _GEN_3596; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3598 = 12'he0e == io_in ? 12'hed1 : _GEN_3597; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3599 = 12'he0f == io_in ? 12'hd6b : _GEN_3598; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3600 = 12'he10 == io_in ? 12'ha66 : _GEN_3599; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3601 = 12'he11 == io_in ? 12'hcca : _GEN_3600; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3602 = 12'he12 == io_in ? 12'hf2f : _GEN_3601; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3603 = 12'he13 == io_in ? 12'h1e1 : _GEN_3602; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3604 = 12'he14 == io_in ? 12'h1c3 : _GEN_3603; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3605 = 12'he15 == io_in ? 12'hdb9 : _GEN_3604; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3606 = 12'he16 == io_in ? 12'h5d9 : _GEN_3605; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3607 = 12'he17 == io_in ? 12'h254 : _GEN_3606; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3608 = 12'he18 == io_in ? 12'hcae : _GEN_3607; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3609 = 12'he19 == io_in ? 12'hbb6 : _GEN_3608; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3610 = 12'he1a == io_in ? 12'hde7 : _GEN_3609; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3611 = 12'he1b == io_in ? 12'hade : _GEN_3610; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3612 = 12'he1c == io_in ? 12'h24f : _GEN_3611; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3613 = 12'he1d == io_in ? 12'h6b : _GEN_3612; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3614 = 12'he1e == io_in ? 12'hd11 : _GEN_3613; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3615 = 12'he1f == io_in ? 12'h653 : _GEN_3614; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3616 = 12'he20 == io_in ? 12'h1c0 : _GEN_3615; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3617 = 12'he21 == io_in ? 12'hb42 : _GEN_3616; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3618 = 12'he22 == io_in ? 12'h1d9 : _GEN_3617; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3619 = 12'he23 == io_in ? 12'h487 : _GEN_3618; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3620 = 12'he24 == io_in ? 12'hf1e : _GEN_3619; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3621 = 12'he25 == io_in ? 12'ha76 : _GEN_3620; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3622 = 12'he26 == io_in ? 12'h623 : _GEN_3621; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3623 = 12'he27 == io_in ? 12'h90 : _GEN_3622; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3624 = 12'he28 == io_in ? 12'h687 : _GEN_3623; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3625 = 12'he29 == io_in ? 12'h8e2 : _GEN_3624; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3626 = 12'he2a == io_in ? 12'hb7c : _GEN_3625; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3627 = 12'he2b == io_in ? 12'h382 : _GEN_3626; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3628 = 12'he2c == io_in ? 12'h6fd : _GEN_3627; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3629 = 12'he2d == io_in ? 12'ha9b : _GEN_3628; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3630 = 12'he2e == io_in ? 12'h880 : _GEN_3629; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3631 = 12'he2f == io_in ? 12'h42f : _GEN_3630; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3632 = 12'he30 == io_in ? 12'h8e7 : _GEN_3631; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3633 = 12'he31 == io_in ? 12'ha5e : _GEN_3632; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3634 = 12'he32 == io_in ? 12'haa3 : _GEN_3633; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3635 = 12'he33 == io_in ? 12'h13e : _GEN_3634; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3636 = 12'he34 == io_in ? 12'h549 : _GEN_3635; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3637 = 12'he35 == io_in ? 12'h7b9 : _GEN_3636; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3638 = 12'he36 == io_in ? 12'h897 : _GEN_3637; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3639 = 12'he37 == io_in ? 12'h657 : _GEN_3638; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3640 = 12'he38 == io_in ? 12'h350 : _GEN_3639; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3641 = 12'he39 == io_in ? 12'h150 : _GEN_3640; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3642 = 12'he3a == io_in ? 12'h6a : _GEN_3641; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3643 = 12'he3b == io_in ? 12'h15c : _GEN_3642; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3644 = 12'he3c == io_in ? 12'h82d : _GEN_3643; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3645 = 12'he3d == io_in ? 12'hd62 : _GEN_3644; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3646 = 12'he3e == io_in ? 12'h362 : _GEN_3645; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3647 = 12'he3f == io_in ? 12'hc96 : _GEN_3646; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3648 = 12'he40 == io_in ? 12'h449 : _GEN_3647; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3649 = 12'he41 == io_in ? 12'hd0f : _GEN_3648; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3650 = 12'he42 == io_in ? 12'hff5 : _GEN_3649; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3651 = 12'he43 == io_in ? 12'hc85 : _GEN_3650; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3652 = 12'he44 == io_in ? 12'h14c : _GEN_3651; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3653 = 12'he45 == io_in ? 12'hb28 : _GEN_3652; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3654 = 12'he46 == io_in ? 12'h70 : _GEN_3653; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3655 = 12'he47 == io_in ? 12'hb57 : _GEN_3654; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3656 = 12'he48 == io_in ? 12'hb89 : _GEN_3655; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3657 = 12'he49 == io_in ? 12'he2d : _GEN_3656; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3658 = 12'he4a == io_in ? 12'h8de : _GEN_3657; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3659 = 12'he4b == io_in ? 12'hba6 : _GEN_3658; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3660 = 12'he4c == io_in ? 12'h2cd : _GEN_3659; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3661 = 12'he4d == io_in ? 12'hd5e : _GEN_3660; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3662 = 12'he4e == io_in ? 12'hfad : _GEN_3661; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3663 = 12'he4f == io_in ? 12'h3c2 : _GEN_3662; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3664 = 12'he50 == io_in ? 12'h1a3 : _GEN_3663; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3665 = 12'he51 == io_in ? 12'hbcf : _GEN_3664; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3666 = 12'he52 == io_in ? 12'h683 : _GEN_3665; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3667 = 12'he53 == io_in ? 12'ha56 : _GEN_3666; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3668 = 12'he54 == io_in ? 12'h530 : _GEN_3667; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3669 = 12'he55 == io_in ? 12'h131 : _GEN_3668; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3670 = 12'he56 == io_in ? 12'h99d : _GEN_3669; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3671 = 12'he57 == io_in ? 12'h44f : _GEN_3670; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3672 = 12'he58 == io_in ? 12'hcb9 : _GEN_3671; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3673 = 12'he59 == io_in ? 12'h8ab : _GEN_3672; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3674 = 12'he5a == io_in ? 12'h63f : _GEN_3673; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3675 = 12'he5b == io_in ? 12'h756 : _GEN_3674; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3676 = 12'he5c == io_in ? 12'h757 : _GEN_3675; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3677 = 12'he5d == io_in ? 12'ha18 : _GEN_3676; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3678 = 12'he5e == io_in ? 12'h90e : _GEN_3677; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3679 = 12'he5f == io_in ? 12'hfd9 : _GEN_3678; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3680 = 12'he60 == io_in ? 12'h51e : _GEN_3679; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3681 = 12'he61 == io_in ? 12'h3cc : _GEN_3680; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3682 = 12'he62 == io_in ? 12'h3e7 : _GEN_3681; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3683 = 12'he63 == io_in ? 12'hefb : _GEN_3682; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3684 = 12'he64 == io_in ? 12'h98a : _GEN_3683; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3685 = 12'he65 == io_in ? 12'hac8 : _GEN_3684; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3686 = 12'he66 == io_in ? 12'h39b : _GEN_3685; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3687 = 12'he67 == io_in ? 12'hc0c : _GEN_3686; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3688 = 12'he68 == io_in ? 12'hf4e : _GEN_3687; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3689 = 12'he69 == io_in ? 12'hfae : _GEN_3688; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3690 = 12'he6a == io_in ? 12'hfc4 : _GEN_3689; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3691 = 12'he6b == io_in ? 12'h484 : _GEN_3690; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3692 = 12'he6c == io_in ? 12'he4e : _GEN_3691; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3693 = 12'he6d == io_in ? 12'h8f4 : _GEN_3692; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3694 = 12'he6e == io_in ? 12'h394 : _GEN_3693; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3695 = 12'he6f == io_in ? 12'h182 : _GEN_3694; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3696 = 12'he70 == io_in ? 12'h603 : _GEN_3695; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3697 = 12'he71 == io_in ? 12'h992 : _GEN_3696; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3698 = 12'he72 == io_in ? 12'hb7a : _GEN_3697; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3699 = 12'he73 == io_in ? 12'hd25 : _GEN_3698; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3700 = 12'he74 == io_in ? 12'h40 : _GEN_3699; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3701 = 12'he75 == io_in ? 12'h4c : _GEN_3700; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3702 = 12'he76 == io_in ? 12'h16e : _GEN_3701; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3703 = 12'he77 == io_in ? 12'hdf2 : _GEN_3702; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3704 = 12'he78 == io_in ? 12'h6b7 : _GEN_3703; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3705 = 12'he79 == io_in ? 12'ha75 : _GEN_3704; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3706 = 12'he7a == io_in ? 12'hc47 : _GEN_3705; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3707 = 12'he7b == io_in ? 12'h1dd : _GEN_3706; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3708 = 12'he7c == io_in ? 12'hb25 : _GEN_3707; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3709 = 12'he7d == io_in ? 12'hf4b : _GEN_3708; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3710 = 12'he7e == io_in ? 12'h4dd : _GEN_3709; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3711 = 12'he7f == io_in ? 12'hb4b : _GEN_3710; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3712 = 12'he80 == io_in ? 12'hd49 : _GEN_3711; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3713 = 12'he81 == io_in ? 12'hb3d : _GEN_3712; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3714 = 12'he82 == io_in ? 12'h83e : _GEN_3713; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3715 = 12'he83 == io_in ? 12'h3e1 : _GEN_3714; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3716 = 12'he84 == io_in ? 12'hfe4 : _GEN_3715; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3717 = 12'he85 == io_in ? 12'h699 : _GEN_3716; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3718 = 12'he86 == io_in ? 12'he73 : _GEN_3717; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3719 = 12'he87 == io_in ? 12'hda7 : _GEN_3718; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3720 = 12'he88 == io_in ? 12'h7fa : _GEN_3719; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3721 = 12'he89 == io_in ? 12'h660 : _GEN_3720; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3722 = 12'he8a == io_in ? 12'h1fc : _GEN_3721; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3723 = 12'he8b == io_in ? 12'habb : _GEN_3722; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3724 = 12'he8c == io_in ? 12'hee4 : _GEN_3723; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3725 = 12'he8d == io_in ? 12'hac0 : _GEN_3724; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3726 = 12'he8e == io_in ? 12'h18a : _GEN_3725; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3727 = 12'he8f == io_in ? 12'h578 : _GEN_3726; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3728 = 12'he90 == io_in ? 12'hc55 : _GEN_3727; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3729 = 12'he91 == io_in ? 12'h255 : _GEN_3728; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3730 = 12'he92 == io_in ? 12'haac : _GEN_3729; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3731 = 12'he93 == io_in ? 12'h2f2 : _GEN_3730; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3732 = 12'he94 == io_in ? 12'h2fb : _GEN_3731; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3733 = 12'he95 == io_in ? 12'h762 : _GEN_3732; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3734 = 12'he96 == io_in ? 12'hbf0 : _GEN_3733; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3735 = 12'he97 == io_in ? 12'hb64 : _GEN_3734; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3736 = 12'he98 == io_in ? 12'h730 : _GEN_3735; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3737 = 12'he99 == io_in ? 12'h1de : _GEN_3736; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3738 = 12'he9a == io_in ? 12'hd03 : _GEN_3737; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3739 = 12'he9b == io_in ? 12'h865 : _GEN_3738; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3740 = 12'he9c == io_in ? 12'hfd7 : _GEN_3739; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3741 = 12'he9d == io_in ? 12'hadc : _GEN_3740; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3742 = 12'he9e == io_in ? 12'hcd8 : _GEN_3741; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3743 = 12'he9f == io_in ? 12'hfbd : _GEN_3742; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3744 = 12'hea0 == io_in ? 12'h639 : _GEN_3743; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3745 = 12'hea1 == io_in ? 12'h94b : _GEN_3744; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3746 = 12'hea2 == io_in ? 12'h52e : _GEN_3745; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3747 = 12'hea3 == io_in ? 12'h26 : _GEN_3746; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3748 = 12'hea4 == io_in ? 12'ha66 : _GEN_3747; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3749 = 12'hea5 == io_in ? 12'h1d9 : _GEN_3748; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3750 = 12'hea6 == io_in ? 12'hf23 : _GEN_3749; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3751 = 12'hea7 == io_in ? 12'h886 : _GEN_3750; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3752 = 12'hea8 == io_in ? 12'h20 : _GEN_3751; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3753 = 12'hea9 == io_in ? 12'ha85 : _GEN_3752; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3754 = 12'heaa == io_in ? 12'h185 : _GEN_3753; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3755 = 12'heab == io_in ? 12'h31a : _GEN_3754; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3756 = 12'heac == io_in ? 12'hf99 : _GEN_3755; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3757 = 12'head == io_in ? 12'h309 : _GEN_3756; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3758 = 12'heae == io_in ? 12'hc24 : _GEN_3757; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3759 = 12'heaf == io_in ? 12'h687 : _GEN_3758; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3760 = 12'heb0 == io_in ? 12'h9c2 : _GEN_3759; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3761 = 12'heb1 == io_in ? 12'hcc1 : _GEN_3760; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3762 = 12'heb2 == io_in ? 12'h620 : _GEN_3761; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3763 = 12'heb3 == io_in ? 12'hc2e : _GEN_3762; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3764 = 12'heb4 == io_in ? 12'h662 : _GEN_3763; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3765 = 12'heb5 == io_in ? 12'hcbc : _GEN_3764; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3766 = 12'heb6 == io_in ? 12'hbac : _GEN_3765; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3767 = 12'heb7 == io_in ? 12'h3e9 : _GEN_3766; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3768 = 12'heb8 == io_in ? 12'h24d : _GEN_3767; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3769 = 12'heb9 == io_in ? 12'h882 : _GEN_3768; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3770 = 12'heba == io_in ? 12'h249 : _GEN_3769; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3771 = 12'hebb == io_in ? 12'h363 : _GEN_3770; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3772 = 12'hebc == io_in ? 12'hcc9 : _GEN_3771; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3773 = 12'hebd == io_in ? 12'hff2 : _GEN_3772; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3774 = 12'hebe == io_in ? 12'h423 : _GEN_3773; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3775 = 12'hebf == io_in ? 12'h554 : _GEN_3774; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3776 = 12'hec0 == io_in ? 12'hea2 : _GEN_3775; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3777 = 12'hec1 == io_in ? 12'h492 : _GEN_3776; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3778 = 12'hec2 == io_in ? 12'h21e : _GEN_3777; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3779 = 12'hec3 == io_in ? 12'h997 : _GEN_3778; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3780 = 12'hec4 == io_in ? 12'hd49 : _GEN_3779; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3781 = 12'hec5 == io_in ? 12'h6d2 : _GEN_3780; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3782 = 12'hec6 == io_in ? 12'ha16 : _GEN_3781; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3783 = 12'hec7 == io_in ? 12'h9a4 : _GEN_3782; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3784 = 12'hec8 == io_in ? 12'hcd9 : _GEN_3783; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3785 = 12'hec9 == io_in ? 12'h54f : _GEN_3784; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3786 = 12'heca == io_in ? 12'h874 : _GEN_3785; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3787 = 12'hecb == io_in ? 12'h84c : _GEN_3786; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3788 = 12'hecc == io_in ? 12'h1bc : _GEN_3787; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3789 = 12'hecd == io_in ? 12'hf66 : _GEN_3788; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3790 = 12'hece == io_in ? 12'h9b9 : _GEN_3789; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3791 = 12'hecf == io_in ? 12'h3ac : _GEN_3790; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3792 = 12'hed0 == io_in ? 12'hc13 : _GEN_3791; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3793 = 12'hed1 == io_in ? 12'h4ca : _GEN_3792; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3794 = 12'hed2 == io_in ? 12'h577 : _GEN_3793; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3795 = 12'hed3 == io_in ? 12'hc62 : _GEN_3794; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3796 = 12'hed4 == io_in ? 12'hb83 : _GEN_3795; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3797 = 12'hed5 == io_in ? 12'h6ea : _GEN_3796; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3798 = 12'hed6 == io_in ? 12'he5e : _GEN_3797; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3799 = 12'hed7 == io_in ? 12'h5a8 : _GEN_3798; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3800 = 12'hed8 == io_in ? 12'ha71 : _GEN_3799; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3801 = 12'hed9 == io_in ? 12'hfdc : _GEN_3800; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3802 = 12'heda == io_in ? 12'hd58 : _GEN_3801; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3803 = 12'hedb == io_in ? 12'hb06 : _GEN_3802; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3804 = 12'hedc == io_in ? 12'h57a : _GEN_3803; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3805 = 12'hedd == io_in ? 12'hdb7 : _GEN_3804; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3806 = 12'hede == io_in ? 12'h41b : _GEN_3805; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3807 = 12'hedf == io_in ? 12'he55 : _GEN_3806; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3808 = 12'hee0 == io_in ? 12'h32c : _GEN_3807; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3809 = 12'hee1 == io_in ? 12'ha79 : _GEN_3808; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3810 = 12'hee2 == io_in ? 12'h78b : _GEN_3809; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3811 = 12'hee3 == io_in ? 12'hcd8 : _GEN_3810; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3812 = 12'hee4 == io_in ? 12'hbe7 : _GEN_3811; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3813 = 12'hee5 == io_in ? 12'h70 : _GEN_3812; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3814 = 12'hee6 == io_in ? 12'h634 : _GEN_3813; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3815 = 12'hee7 == io_in ? 12'hce5 : _GEN_3814; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3816 = 12'hee8 == io_in ? 12'h1a7 : _GEN_3815; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3817 = 12'hee9 == io_in ? 12'h423 : _GEN_3816; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3818 = 12'heea == io_in ? 12'hb23 : _GEN_3817; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3819 = 12'heeb == io_in ? 12'hc91 : _GEN_3818; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3820 = 12'heec == io_in ? 12'h853 : _GEN_3819; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3821 = 12'heed == io_in ? 12'hfc3 : _GEN_3820; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3822 = 12'heee == io_in ? 12'h22e : _GEN_3821; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3823 = 12'heef == io_in ? 12'h247 : _GEN_3822; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3824 = 12'hef0 == io_in ? 12'hb4e : _GEN_3823; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3825 = 12'hef1 == io_in ? 12'hc94 : _GEN_3824; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3826 = 12'hef2 == io_in ? 12'hef4 : _GEN_3825; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3827 = 12'hef3 == io_in ? 12'hc2c : _GEN_3826; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3828 = 12'hef4 == io_in ? 12'hbdb : _GEN_3827; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3829 = 12'hef5 == io_in ? 12'h5a2 : _GEN_3828; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3830 = 12'hef6 == io_in ? 12'hadb : _GEN_3829; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3831 = 12'hef7 == io_in ? 12'h478 : _GEN_3830; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3832 = 12'hef8 == io_in ? 12'h205 : _GEN_3831; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3833 = 12'hef9 == io_in ? 12'h4c : _GEN_3832; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3834 = 12'hefa == io_in ? 12'hd2b : _GEN_3833; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3835 = 12'hefb == io_in ? 12'hdf2 : _GEN_3834; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3836 = 12'hefc == io_in ? 12'h962 : _GEN_3835; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3837 = 12'hefd == io_in ? 12'h49b : _GEN_3836; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3838 = 12'hefe == io_in ? 12'h8d4 : _GEN_3837; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3839 = 12'heff == io_in ? 12'h2f4 : _GEN_3838; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3840 = 12'hf00 == io_in ? 12'h2ef : _GEN_3839; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3841 = 12'hf01 == io_in ? 12'hcdc : _GEN_3840; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3842 = 12'hf02 == io_in ? 12'h934 : _GEN_3841; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3843 = 12'hf03 == io_in ? 12'hd69 : _GEN_3842; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3844 = 12'hf04 == io_in ? 12'h28a : _GEN_3843; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3845 = 12'hf05 == io_in ? 12'h473 : _GEN_3844; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3846 = 12'hf06 == io_in ? 12'h668 : _GEN_3845; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3847 = 12'hf07 == io_in ? 12'h26f : _GEN_3846; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3848 = 12'hf08 == io_in ? 12'ha23 : _GEN_3847; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3849 = 12'hf09 == io_in ? 12'h563 : _GEN_3848; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3850 = 12'hf0a == io_in ? 12'hcbb : _GEN_3849; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3851 = 12'hf0b == io_in ? 12'h78b : _GEN_3850; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3852 = 12'hf0c == io_in ? 12'h64e : _GEN_3851; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3853 = 12'hf0d == io_in ? 12'hded : _GEN_3852; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3854 = 12'hf0e == io_in ? 12'h415 : _GEN_3853; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3855 = 12'hf0f == io_in ? 12'h97a : _GEN_3854; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3856 = 12'hf10 == io_in ? 12'hb13 : _GEN_3855; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3857 = 12'hf11 == io_in ? 12'h8e4 : _GEN_3856; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3858 = 12'hf12 == io_in ? 12'hcd2 : _GEN_3857; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3859 = 12'hf13 == io_in ? 12'h955 : _GEN_3858; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3860 = 12'hf14 == io_in ? 12'h683 : _GEN_3859; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3861 = 12'hf15 == io_in ? 12'hf39 : _GEN_3860; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3862 = 12'hf16 == io_in ? 12'h3c : _GEN_3861; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3863 = 12'hf17 == io_in ? 12'h7c6 : _GEN_3862; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3864 = 12'hf18 == io_in ? 12'h716 : _GEN_3863; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3865 = 12'hf19 == io_in ? 12'h5b0 : _GEN_3864; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3866 = 12'hf1a == io_in ? 12'hb2a : _GEN_3865; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3867 = 12'hf1b == io_in ? 12'h81d : _GEN_3866; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3868 = 12'hf1c == io_in ? 12'ha90 : _GEN_3867; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3869 = 12'hf1d == io_in ? 12'h232 : _GEN_3868; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3870 = 12'hf1e == io_in ? 12'h8d9 : _GEN_3869; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3871 = 12'hf1f == io_in ? 12'he3d : _GEN_3870; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3872 = 12'hf20 == io_in ? 12'h7c4 : _GEN_3871; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3873 = 12'hf21 == io_in ? 12'hf49 : _GEN_3872; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3874 = 12'hf22 == io_in ? 12'h9b : _GEN_3873; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3875 = 12'hf23 == io_in ? 12'h7bf : _GEN_3874; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3876 = 12'hf24 == io_in ? 12'hff : _GEN_3875; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3877 = 12'hf25 == io_in ? 12'h627 : _GEN_3876; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3878 = 12'hf26 == io_in ? 12'h87d : _GEN_3877; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3879 = 12'hf27 == io_in ? 12'h711 : _GEN_3878; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3880 = 12'hf28 == io_in ? 12'h185 : _GEN_3879; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3881 = 12'hf29 == io_in ? 12'h6cf : _GEN_3880; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3882 = 12'hf2a == io_in ? 12'he04 : _GEN_3881; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3883 = 12'hf2b == io_in ? 12'h817 : _GEN_3882; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3884 = 12'hf2c == io_in ? 12'h79b : _GEN_3883; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3885 = 12'hf2d == io_in ? 12'hfb6 : _GEN_3884; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3886 = 12'hf2e == io_in ? 12'h918 : _GEN_3885; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3887 = 12'hf2f == io_in ? 12'h295 : _GEN_3886; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3888 = 12'hf30 == io_in ? 12'h3db : _GEN_3887; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3889 = 12'hf31 == io_in ? 12'h122 : _GEN_3888; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3890 = 12'hf32 == io_in ? 12'h6ee : _GEN_3889; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3891 = 12'hf33 == io_in ? 12'hce7 : _GEN_3890; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3892 = 12'hf34 == io_in ? 12'h236 : _GEN_3891; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3893 = 12'hf35 == io_in ? 12'haa7 : _GEN_3892; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3894 = 12'hf36 == io_in ? 12'he68 : _GEN_3893; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3895 = 12'hf37 == io_in ? 12'hf82 : _GEN_3894; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3896 = 12'hf38 == io_in ? 12'hba : _GEN_3895; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3897 = 12'hf39 == io_in ? 12'h186 : _GEN_3896; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3898 = 12'hf3a == io_in ? 12'h625 : _GEN_3897; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3899 = 12'hf3b == io_in ? 12'h1a9 : _GEN_3898; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3900 = 12'hf3c == io_in ? 12'h326 : _GEN_3899; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3901 = 12'hf3d == io_in ? 12'hb95 : _GEN_3900; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3902 = 12'hf3e == io_in ? 12'h42 : _GEN_3901; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3903 = 12'hf3f == io_in ? 12'h405 : _GEN_3902; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3904 = 12'hf40 == io_in ? 12'ha64 : _GEN_3903; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3905 = 12'hf41 == io_in ? 12'hbc6 : _GEN_3904; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3906 = 12'hf42 == io_in ? 12'hfd4 : _GEN_3905; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3907 = 12'hf43 == io_in ? 12'hd6a : _GEN_3906; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3908 = 12'hf44 == io_in ? 12'he00 : _GEN_3907; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3909 = 12'hf45 == io_in ? 12'h9b1 : _GEN_3908; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3910 = 12'hf46 == io_in ? 12'h146 : _GEN_3909; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3911 = 12'hf47 == io_in ? 12'h7be : _GEN_3910; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3912 = 12'hf48 == io_in ? 12'hff4 : _GEN_3911; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3913 = 12'hf49 == io_in ? 12'hd73 : _GEN_3912; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3914 = 12'hf4a == io_in ? 12'he87 : _GEN_3913; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3915 = 12'hf4b == io_in ? 12'h23c : _GEN_3914; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3916 = 12'hf4c == io_in ? 12'hcff : _GEN_3915; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3917 = 12'hf4d == io_in ? 12'hba1 : _GEN_3916; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3918 = 12'hf4e == io_in ? 12'h1b8 : _GEN_3917; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3919 = 12'hf4f == io_in ? 12'h697 : _GEN_3918; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3920 = 12'hf50 == io_in ? 12'hbfa : _GEN_3919; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3921 = 12'hf51 == io_in ? 12'haeb : _GEN_3920; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3922 = 12'hf52 == io_in ? 12'h8bd : _GEN_3921; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3923 = 12'hf53 == io_in ? 12'hf65 : _GEN_3922; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3924 = 12'hf54 == io_in ? 12'hc1c : _GEN_3923; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3925 = 12'hf55 == io_in ? 12'he16 : _GEN_3924; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3926 = 12'hf56 == io_in ? 12'hfdc : _GEN_3925; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3927 = 12'hf57 == io_in ? 12'h824 : _GEN_3926; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3928 = 12'hf58 == io_in ? 12'h651 : _GEN_3927; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3929 = 12'hf59 == io_in ? 12'haa4 : _GEN_3928; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3930 = 12'hf5a == io_in ? 12'h39e : _GEN_3929; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3931 = 12'hf5b == io_in ? 12'hddd : _GEN_3930; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3932 = 12'hf5c == io_in ? 12'h19a : _GEN_3931; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3933 = 12'hf5d == io_in ? 12'he62 : _GEN_3932; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3934 = 12'hf5e == io_in ? 12'h71e : _GEN_3933; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3935 = 12'hf5f == io_in ? 12'h7f3 : _GEN_3934; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3936 = 12'hf60 == io_in ? 12'ha56 : _GEN_3935; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3937 = 12'hf61 == io_in ? 12'h730 : _GEN_3936; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3938 = 12'hf62 == io_in ? 12'h4a8 : _GEN_3937; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3939 = 12'hf63 == io_in ? 12'h34b : _GEN_3938; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3940 = 12'hf64 == io_in ? 12'hb6d : _GEN_3939; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3941 = 12'hf65 == io_in ? 12'hfec : _GEN_3940; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3942 = 12'hf66 == io_in ? 12'he17 : _GEN_3941; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3943 = 12'hf67 == io_in ? 12'h813 : _GEN_3942; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3944 = 12'hf68 == io_in ? 12'h5a7 : _GEN_3943; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3945 = 12'hf69 == io_in ? 12'hf22 : _GEN_3944; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3946 = 12'hf6a == io_in ? 12'h807 : _GEN_3945; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3947 = 12'hf6b == io_in ? 12'h122 : _GEN_3946; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3948 = 12'hf6c == io_in ? 12'h2c6 : _GEN_3947; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3949 = 12'hf6d == io_in ? 12'h825 : _GEN_3948; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3950 = 12'hf6e == io_in ? 12'h5d : _GEN_3949; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3951 = 12'hf6f == io_in ? 12'hb5 : _GEN_3950; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3952 = 12'hf70 == io_in ? 12'h879 : _GEN_3951; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3953 = 12'hf71 == io_in ? 12'h932 : _GEN_3952; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3954 = 12'hf72 == io_in ? 12'hb95 : _GEN_3953; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3955 = 12'hf73 == io_in ? 12'h304 : _GEN_3954; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3956 = 12'hf74 == io_in ? 12'hb71 : _GEN_3955; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3957 = 12'hf75 == io_in ? 12'ha0d : _GEN_3956; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3958 = 12'hf76 == io_in ? 12'hcd5 : _GEN_3957; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3959 = 12'hf77 == io_in ? 12'h5b8 : _GEN_3958; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3960 = 12'hf78 == io_in ? 12'h889 : _GEN_3959; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3961 = 12'hf79 == io_in ? 12'h281 : _GEN_3960; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3962 = 12'hf7a == io_in ? 12'hf67 : _GEN_3961; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3963 = 12'hf7b == io_in ? 12'h225 : _GEN_3962; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3964 = 12'hf7c == io_in ? 12'h3ca : _GEN_3963; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3965 = 12'hf7d == io_in ? 12'h3e : _GEN_3964; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3966 = 12'hf7e == io_in ? 12'hb24 : _GEN_3965; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3967 = 12'hf7f == io_in ? 12'hd95 : _GEN_3966; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3968 = 12'hf80 == io_in ? 12'h1ac : _GEN_3967; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3969 = 12'hf81 == io_in ? 12'hd1f : _GEN_3968; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3970 = 12'hf82 == io_in ? 12'h400 : _GEN_3969; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3971 = 12'hf83 == io_in ? 12'h9e0 : _GEN_3970; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3972 = 12'hf84 == io_in ? 12'h357 : _GEN_3971; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3973 = 12'hf85 == io_in ? 12'h2d6 : _GEN_3972; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3974 = 12'hf86 == io_in ? 12'h390 : _GEN_3973; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3975 = 12'hf87 == io_in ? 12'h3f7 : _GEN_3974; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3976 = 12'hf88 == io_in ? 12'hbdc : _GEN_3975; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3977 = 12'hf89 == io_in ? 12'h588 : _GEN_3976; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3978 = 12'hf8a == io_in ? 12'hc3e : _GEN_3977; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3979 = 12'hf8b == io_in ? 12'h51e : _GEN_3978; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3980 = 12'hf8c == io_in ? 12'ha3b : _GEN_3979; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3981 = 12'hf8d == io_in ? 12'hd7d : _GEN_3980; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3982 = 12'hf8e == io_in ? 12'hbb0 : _GEN_3981; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3983 = 12'hf8f == io_in ? 12'hdfb : _GEN_3982; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3984 = 12'hf90 == io_in ? 12'hdb8 : _GEN_3983; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3985 = 12'hf91 == io_in ? 12'h6f5 : _GEN_3984; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3986 = 12'hf92 == io_in ? 12'hd43 : _GEN_3985; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3987 = 12'hf93 == io_in ? 12'hbfb : _GEN_3986; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3988 = 12'hf94 == io_in ? 12'h1f0 : _GEN_3987; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3989 = 12'hf95 == io_in ? 12'h91f : _GEN_3988; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3990 = 12'hf96 == io_in ? 12'hfbf : _GEN_3989; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3991 = 12'hf97 == io_in ? 12'he04 : _GEN_3990; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3992 = 12'hf98 == io_in ? 12'h43e : _GEN_3991; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3993 = 12'hf99 == io_in ? 12'h805 : _GEN_3992; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3994 = 12'hf9a == io_in ? 12'h189 : _GEN_3993; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3995 = 12'hf9b == io_in ? 12'hd29 : _GEN_3994; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3996 = 12'hf9c == io_in ? 12'h8e2 : _GEN_3995; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3997 = 12'hf9d == io_in ? 12'h4f1 : _GEN_3996; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3998 = 12'hf9e == io_in ? 12'h4b9 : _GEN_3997; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_3999 = 12'hf9f == io_in ? 12'h982 : _GEN_3998; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4000 = 12'hfa0 == io_in ? 12'hc94 : _GEN_3999; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4001 = 12'hfa1 == io_in ? 12'hb66 : _GEN_4000; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4002 = 12'hfa2 == io_in ? 12'h5a6 : _GEN_4001; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4003 = 12'hfa3 == io_in ? 12'h793 : _GEN_4002; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4004 = 12'hfa4 == io_in ? 12'h5d5 : _GEN_4003; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4005 = 12'hfa5 == io_in ? 12'ha8a : _GEN_4004; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4006 = 12'hfa6 == io_in ? 12'h1b8 : _GEN_4005; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4007 = 12'hfa7 == io_in ? 12'h43a : _GEN_4006; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4008 = 12'hfa8 == io_in ? 12'h397 : _GEN_4007; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4009 = 12'hfa9 == io_in ? 12'h2c7 : _GEN_4008; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4010 = 12'hfaa == io_in ? 12'hcf6 : _GEN_4009; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4011 = 12'hfab == io_in ? 12'h5d1 : _GEN_4010; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4012 = 12'hfac == io_in ? 12'hdf9 : _GEN_4011; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4013 = 12'hfad == io_in ? 12'h205 : _GEN_4012; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4014 = 12'hfae == io_in ? 12'h48 : _GEN_4013; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4015 = 12'hfaf == io_in ? 12'h1fb : _GEN_4014; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4016 = 12'hfb0 == io_in ? 12'h7e9 : _GEN_4015; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4017 = 12'hfb1 == io_in ? 12'h57e : _GEN_4016; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4018 = 12'hfb2 == io_in ? 12'haf2 : _GEN_4017; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4019 = 12'hfb3 == io_in ? 12'hee5 : _GEN_4018; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4020 = 12'hfb4 == io_in ? 12'h115 : _GEN_4019; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4021 = 12'hfb5 == io_in ? 12'hc32 : _GEN_4020; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4022 = 12'hfb6 == io_in ? 12'h2f2 : _GEN_4021; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4023 = 12'hfb7 == io_in ? 12'h9b7 : _GEN_4022; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4024 = 12'hfb8 == io_in ? 12'h720 : _GEN_4023; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4025 = 12'hfb9 == io_in ? 12'hff5 : _GEN_4024; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4026 = 12'hfba == io_in ? 12'h287 : _GEN_4025; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4027 = 12'hfbb == io_in ? 12'h5ea : _GEN_4026; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4028 = 12'hfbc == io_in ? 12'h213 : _GEN_4027; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4029 = 12'hfbd == io_in ? 12'h309 : _GEN_4028; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4030 = 12'hfbe == io_in ? 12'hf49 : _GEN_4029; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4031 = 12'hfbf == io_in ? 12'hb92 : _GEN_4030; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4032 = 12'hfc0 == io_in ? 12'hcb4 : _GEN_4031; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4033 = 12'hfc1 == io_in ? 12'h519 : _GEN_4032; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4034 = 12'hfc2 == io_in ? 12'h856 : _GEN_4033; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4035 = 12'hfc3 == io_in ? 12'hd29 : _GEN_4034; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4036 = 12'hfc4 == io_in ? 12'hfae : _GEN_4035; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4037 = 12'hfc5 == io_in ? 12'h2cc : _GEN_4036; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4038 = 12'hfc6 == io_in ? 12'h562 : _GEN_4037; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4039 = 12'hfc7 == io_in ? 12'he5a : _GEN_4038; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4040 = 12'hfc8 == io_in ? 12'ha35 : _GEN_4039; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4041 = 12'hfc9 == io_in ? 12'hfa3 : _GEN_4040; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4042 = 12'hfca == io_in ? 12'h66a : _GEN_4041; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4043 = 12'hfcb == io_in ? 12'h4c : _GEN_4042; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4044 = 12'hfcc == io_in ? 12'h904 : _GEN_4043; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4045 = 12'hfcd == io_in ? 12'h92f : _GEN_4044; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4046 = 12'hfce == io_in ? 12'h9ae : _GEN_4045; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4047 = 12'hfcf == io_in ? 12'h885 : _GEN_4046; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4048 = 12'hfd0 == io_in ? 12'h355 : _GEN_4047; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4049 = 12'hfd1 == io_in ? 12'h633 : _GEN_4048; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4050 = 12'hfd2 == io_in ? 12'h867 : _GEN_4049; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4051 = 12'hfd3 == io_in ? 12'hd2e : _GEN_4050; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4052 = 12'hfd4 == io_in ? 12'hc30 : _GEN_4051; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4053 = 12'hfd5 == io_in ? 12'hb50 : _GEN_4052; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4054 = 12'hfd6 == io_in ? 12'hfcd : _GEN_4053; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4055 = 12'hfd7 == io_in ? 12'h4ab : _GEN_4054; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4056 = 12'hfd8 == io_in ? 12'he34 : _GEN_4055; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4057 = 12'hfd9 == io_in ? 12'hae5 : _GEN_4056; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4058 = 12'hfda == io_in ? 12'h5e2 : _GEN_4057; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4059 = 12'hfdb == io_in ? 12'hafb : _GEN_4058; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4060 = 12'hfdc == io_in ? 12'ha11 : _GEN_4059; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4061 = 12'hfdd == io_in ? 12'hf1a : _GEN_4060; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4062 = 12'hfde == io_in ? 12'hcea : _GEN_4061; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4063 = 12'hfdf == io_in ? 12'ha21 : _GEN_4062; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4064 = 12'hfe0 == io_in ? 12'h5d : _GEN_4063; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4065 = 12'hfe1 == io_in ? 12'h52a : _GEN_4064; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4066 = 12'hfe2 == io_in ? 12'h61c : _GEN_4065; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4067 = 12'hfe3 == io_in ? 12'hc35 : _GEN_4066; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4068 = 12'hfe4 == io_in ? 12'h1d1 : _GEN_4067; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4069 = 12'hfe5 == io_in ? 12'h928 : _GEN_4068; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4070 = 12'hfe6 == io_in ? 12'heea : _GEN_4069; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4071 = 12'hfe7 == io_in ? 12'h741 : _GEN_4070; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4072 = 12'hfe8 == io_in ? 12'hbd0 : _GEN_4071; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4073 = 12'hfe9 == io_in ? 12'hb44 : _GEN_4072; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4074 = 12'hfea == io_in ? 12'h3fb : _GEN_4073; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4075 = 12'hfeb == io_in ? 12'h953 : _GEN_4074; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4076 = 12'hfec == io_in ? 12'h8b8 : _GEN_4075; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4077 = 12'hfed == io_in ? 12'hd00 : _GEN_4076; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4078 = 12'hfee == io_in ? 12'haa2 : _GEN_4077; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4079 = 12'hfef == io_in ? 12'hc76 : _GEN_4078; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4080 = 12'hff0 == io_in ? 12'hc71 : _GEN_4079; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4081 = 12'hff1 == io_in ? 12'h7fb : _GEN_4080; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4082 = 12'hff2 == io_in ? 12'hb83 : _GEN_4081; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4083 = 12'hff3 == io_in ? 12'h792 : _GEN_4082; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4084 = 12'hff4 == io_in ? 12'hf43 : _GEN_4083; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4085 = 12'hff5 == io_in ? 12'h30f : _GEN_4084; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4086 = 12'hff6 == io_in ? 12'h70d : _GEN_4085; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4087 = 12'hff7 == io_in ? 12'h533 : _GEN_4086; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4088 = 12'hff8 == io_in ? 12'h616 : _GEN_4087; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4089 = 12'hff9 == io_in ? 12'hc3 : _GEN_4088; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4090 = 12'hffa == io_in ? 12'h2f9 : _GEN_4089; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4091 = 12'hffb == io_in ? 12'h9c1 : _GEN_4090; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4092 = 12'hffc == io_in ? 12'hb6e : _GEN_4091; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4093 = 12'hffd == io_in ? 12'h57f : _GEN_4092; // @[RandomLUT.scala 22:{10,10}]
  wire [11:0] _GEN_4094 = 12'hffe == io_in ? 12'hd51 : _GEN_4093; // @[RandomLUT.scala 22:{10,10}]
  assign io_out = 12'hfff == io_in ? 12'h667 : _GEN_4094; // @[RandomLUT.scala 22:{10,10}]
endmodule
module RandomLUTPipe(
  input         clock,
  input         reset,
  input  [11:0] io_in,
  output [11:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [11:0] lut_io_in; // @[RandomLUTPipe.scala 13:19]
  wire [11:0] lut_io_out; // @[RandomLUTPipe.scala 13:19]
  reg [11:0] lut_in; // @[RandomLUTPipe.scala 12:23]
  reg [11:0] lut_out; // @[RandomLUTPipe.scala 15:24]
  RandomLUT lut ( // @[RandomLUTPipe.scala 13:19]
    .io_in(lut_io_in),
    .io_out(lut_io_out)
  );
  assign io_out = lut_out; // @[RandomLUTPipe.scala 17:10]
  assign lut_io_in = lut_in; // @[RandomLUTPipe.scala 14:13]
  always @(posedge clock) begin
    lut_in <= io_in; // @[RandomLUTPipe.scala 12:23]
    lut_out <= lut_io_out; // @[RandomLUTPipe.scala 15:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lut_in = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  lut_out = _RAND_1[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
